`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
turbVZeqJTR6A1zNg2Oz/CPXCBxoL9wXnsjKWOHM+4fvwaQfBZt7fC4WtX030QGY
JzycRUbctEVC1Te7di0DznmGwPtpcFKfGLZfJhYRws0c2N26m2JIXl5NFHwycOdn
j0Rt+ZAFoMtVvW4WbM1GgMkd4xaNsvEjeHCu14/acr9cAR+sb7Y4e0yVgfNESVRI
a3mHIZdLBrzdjawIEnPOFtNjdqafOtzFS29gB+BxMElZ5d/v7nwSd2BmR12KRMhc
xQ0aEkZv7shYkNBSbM2lQHeABT+e/Lu8Sz9fYqnE+DHwVeuTyyCUsGqFlQPCm4am
/FTtMPNx4iycMJmJ7p/AoRlPPnZ4xU3v7AV++O7EyGRE/mY8uvCS2xJgrgdDAk/w
XWa0eXxAjHkZ5eugwB9hy/+GsqXm5tx35ZCac64AlWSgPnuRv2cbw2Rym7N63NWI
ZNvokNbgL3l1BN+WRLZgRJO6h8mr/EXGn0WMLmLIDpAtnkaoxEk9T9kn255IuuUQ
/BP07Xta5Dn9yH2f3z5cqKnMgJ2aRsBII9ygujQzwAr6vCGQxIkbkbM1eXoEwfZ0
+nkHXOOvV80oIt5hZe6iCafjE5DsnfBFKv0Cq6819krtA+UG35mJElmp78DJT9TE
H4weQVHMIX+F+Z60dgx5hfLfpTfHSiOMLjbte46bhCKyFbm3XrlN2sxUh/4qji+q
L2gH69cvTfuKyksQTodK+BTBasyPOyGVmN431nK9qPwfCE5I6SBWecVhOgUB6mjq
qajvJcp77yX0PX7A2VrAwcECkHWcpdGmPMmXOvRwg8kG6RwWX3cJIN2MuXFkYsqa
Hiebt9T8/CQER5nkdJ2VzhBRJDF6D6zFg50XTREuCGTJtTGRZGYTRYQaa4fABQnp
sNhs9WRJElZpfPuyddMHhN/00Bh5T39SYjcBQO4ewc9/tpbBWgBvDOp3Qa+4C1eC
L6M6PriXNi8ovBJ9DzudxrsAcBW8j87t2bS4iPGYtbQ5a41Oul0zvh3vHBOJJS3/
fkGJqv5UF99OnIMCd7fK5IAzjA62t4y0Y4xWFxk3DoQSbe1I0OYrd+uFs2D4JnRR
1vT4939/Nw2x4naSV1a3PvbZa1/ZPd1zwoPXmW3PzZY=
`protect END_PROTECTED
