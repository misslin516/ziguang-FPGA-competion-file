library verilog;
use verilog.vl_types.all;
entity uart_rd_lock is
    port(
        core_clk        : in     vl_logic;
        core_rst_n      : in     vl_logic;
        uart_read_req   : in     vl_logic;
        uart_read_ack   : out    vl_logic;
        uart_read_addr  : in     vl_logic_vector(8 downto 0);
        status_bus_80   : in     vl_logic_vector(31 downto 0);
        status_bus_81   : in     vl_logic_vector(31 downto 0);
        status_bus_82   : in     vl_logic_vector(31 downto 0);
        status_bus_83   : in     vl_logic_vector(31 downto 0);
        status_bus_84   : in     vl_logic_vector(31 downto 0);
        status_bus_85   : in     vl_logic_vector(31 downto 0);
        status_bus_86   : in     vl_logic_vector(31 downto 0);
        status_bus_87   : in     vl_logic_vector(31 downto 0);
        status_bus_88   : in     vl_logic_vector(31 downto 0);
        status_bus_89   : in     vl_logic_vector(31 downto 0);
        status_bus_8a   : in     vl_logic_vector(31 downto 0);
        status_bus_8b   : in     vl_logic_vector(31 downto 0);
        status_bus_8c   : in     vl_logic_vector(31 downto 0);
        status_bus_8d   : in     vl_logic_vector(31 downto 0);
        status_bus_8e   : in     vl_logic_vector(31 downto 0);
        status_bus_8f   : in     vl_logic_vector(31 downto 0);
        status_bus_90   : in     vl_logic_vector(31 downto 0);
        status_bus_91   : in     vl_logic_vector(31 downto 0);
        status_bus_92   : in     vl_logic_vector(31 downto 0);
        status_bus_93   : in     vl_logic_vector(31 downto 0);
        status_bus_94   : in     vl_logic_vector(31 downto 0);
        status_bus_95   : in     vl_logic_vector(31 downto 0);
        status_bus_96   : in     vl_logic_vector(31 downto 0);
        status_bus_97   : in     vl_logic_vector(31 downto 0);
        status_bus_98   : in     vl_logic_vector(31 downto 0);
        status_bus_99   : in     vl_logic_vector(31 downto 0);
        status_bus_9a   : in     vl_logic_vector(31 downto 0);
        status_bus_9b   : in     vl_logic_vector(31 downto 0);
        status_bus_9c   : in     vl_logic_vector(31 downto 0);
        status_bus_9d   : in     vl_logic_vector(31 downto 0);
        status_bus_9e   : in     vl_logic_vector(31 downto 0);
        status_bus_9f   : in     vl_logic_vector(31 downto 0);
        status_bus_a0   : in     vl_logic_vector(31 downto 0);
        status_bus_a1   : in     vl_logic_vector(31 downto 0);
        status_bus_a2   : in     vl_logic_vector(31 downto 0);
        status_bus_a3   : in     vl_logic_vector(31 downto 0);
        status_bus_a4   : in     vl_logic_vector(31 downto 0);
        status_bus_a5   : in     vl_logic_vector(31 downto 0);
        status_bus_a6   : in     vl_logic_vector(31 downto 0);
        status_bus_a7   : in     vl_logic_vector(31 downto 0);
        status_bus_a8   : in     vl_logic_vector(31 downto 0);
        status_bus_a9   : in     vl_logic_vector(31 downto 0);
        status_bus_aa   : in     vl_logic_vector(31 downto 0);
        status_bus_ab   : in     vl_logic_vector(31 downto 0);
        status_bus_ac   : in     vl_logic_vector(31 downto 0);
        status_bus_ad   : in     vl_logic_vector(31 downto 0);
        status_bus_ae   : in     vl_logic_vector(31 downto 0);
        status_bus_af   : in     vl_logic_vector(31 downto 0);
        status_bus_b0   : in     vl_logic_vector(31 downto 0);
        status_bus_b1   : in     vl_logic_vector(31 downto 0);
        status_bus_b2   : in     vl_logic_vector(31 downto 0);
        status_bus_b3   : in     vl_logic_vector(31 downto 0);
        status_bus_b4   : in     vl_logic_vector(31 downto 0);
        status_bus_b5   : in     vl_logic_vector(31 downto 0);
        status_bus_b6   : in     vl_logic_vector(31 downto 0);
        status_bus_b7   : in     vl_logic_vector(31 downto 0);
        status_bus_b8   : in     vl_logic_vector(31 downto 0);
        status_bus_b9   : in     vl_logic_vector(31 downto 0);
        status_bus_ba   : in     vl_logic_vector(31 downto 0);
        status_bus_bb   : in     vl_logic_vector(31 downto 0);
        status_bus_bc   : in     vl_logic_vector(31 downto 0);
        status_bus_bd   : in     vl_logic_vector(31 downto 0);
        status_bus_be   : in     vl_logic_vector(31 downto 0);
        status_bus_bf   : in     vl_logic_vector(31 downto 0);
        status_bus_c0   : in     vl_logic_vector(31 downto 0);
        status_bus_c1   : in     vl_logic_vector(31 downto 0);
        status_bus_c2   : in     vl_logic_vector(31 downto 0);
        status_bus_c3   : in     vl_logic_vector(31 downto 0);
        status_bus_c4   : in     vl_logic_vector(31 downto 0);
        status_bus_c5   : in     vl_logic_vector(31 downto 0);
        status_bus_c6   : in     vl_logic_vector(31 downto 0);
        status_bus_c7   : in     vl_logic_vector(31 downto 0);
        status_bus_c8   : in     vl_logic_vector(31 downto 0);
        status_bus_c9   : in     vl_logic_vector(31 downto 0);
        status_bus_ca   : in     vl_logic_vector(31 downto 0);
        status_bus_cb   : in     vl_logic_vector(31 downto 0);
        status_bus_cc   : in     vl_logic_vector(31 downto 0);
        status_bus_cd   : in     vl_logic_vector(31 downto 0);
        status_bus_ce   : in     vl_logic_vector(31 downto 0);
        status_bus_cf   : in     vl_logic_vector(31 downto 0);
        status_bus_d0   : in     vl_logic_vector(31 downto 0);
        status_bus_d1   : in     vl_logic_vector(31 downto 0);
        status_bus_d2   : in     vl_logic_vector(31 downto 0);
        status_bus_d3   : in     vl_logic_vector(31 downto 0);
        status_bus_d4   : in     vl_logic_vector(31 downto 0);
        status_bus_d5   : in     vl_logic_vector(31 downto 0);
        status_bus_d6   : in     vl_logic_vector(31 downto 0);
        status_bus_d7   : in     vl_logic_vector(31 downto 0);
        status_bus_d8   : in     vl_logic_vector(31 downto 0);
        status_bus_d9   : in     vl_logic_vector(31 downto 0);
        status_bus_da   : in     vl_logic_vector(31 downto 0);
        status_bus_db   : in     vl_logic_vector(31 downto 0);
        status_bus_dc   : in     vl_logic_vector(31 downto 0);
        status_bus_dd   : in     vl_logic_vector(31 downto 0);
        status_bus_de   : in     vl_logic_vector(31 downto 0);
        status_bus_df   : in     vl_logic_vector(31 downto 0);
        status_bus_e0   : in     vl_logic_vector(31 downto 0);
        status_bus_e1   : in     vl_logic_vector(31 downto 0);
        status_bus_e2   : in     vl_logic_vector(31 downto 0);
        status_bus_e3   : in     vl_logic_vector(31 downto 0);
        status_bus_e4   : in     vl_logic_vector(31 downto 0);
        status_bus_e5   : in     vl_logic_vector(31 downto 0);
        status_bus_e6   : in     vl_logic_vector(31 downto 0);
        status_bus_e7   : in     vl_logic_vector(31 downto 0);
        status_bus_e8   : in     vl_logic_vector(31 downto 0);
        status_bus_e9   : in     vl_logic_vector(31 downto 0);
        status_bus_ea   : in     vl_logic_vector(31 downto 0);
        status_bus_eb   : in     vl_logic_vector(31 downto 0);
        status_bus_ec   : in     vl_logic_vector(31 downto 0);
        status_bus_ed   : in     vl_logic_vector(31 downto 0);
        status_bus_ee   : in     vl_logic_vector(31 downto 0);
        status_bus_ef   : in     vl_logic_vector(31 downto 0);
        status_bus_f0   : in     vl_logic_vector(31 downto 0);
        status_bus_f1   : in     vl_logic_vector(31 downto 0);
        status_bus_f2   : in     vl_logic_vector(31 downto 0);
        status_bus_f3   : in     vl_logic_vector(31 downto 0);
        status_bus_f4   : in     vl_logic_vector(31 downto 0);
        status_bus_f5   : in     vl_logic_vector(31 downto 0);
        status_bus_f6   : in     vl_logic_vector(31 downto 0);
        status_bus_f7   : in     vl_logic_vector(31 downto 0);
        status_bus_f8   : in     vl_logic_vector(31 downto 0);
        status_bus_f9   : in     vl_logic_vector(31 downto 0);
        status_bus_fa   : in     vl_logic_vector(31 downto 0);
        status_bus_fb   : in     vl_logic_vector(31 downto 0);
        status_bus_fc   : in     vl_logic_vector(31 downto 0);
        status_bus_fd   : in     vl_logic_vector(31 downto 0);
        status_bus_fe   : in     vl_logic_vector(31 downto 0);
        status_bus_ff   : in     vl_logic_vector(31 downto 0);
        status_bus_lock : out    vl_logic_vector(31 downto 0)
    );
end uart_rd_lock;
