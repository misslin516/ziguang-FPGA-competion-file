`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qj4coVs2R6t3WOVEO0N3YfblogzcA8SkKcBJmbS2g3jY4And35y8tKiMjvz8MkJ
n4iVpfk7gxEITdujnrBe8xwxSyVRqoa6fOQBZyy0J3BiCOBn5LR8/4CNXoNmUotl
cKZPJ0h7IRvHViHufNiN7yuYTjzvvrBLShY/LQTKq7muD7VgxoT+gQVQyCIPXgMd
IoJ+n/LszjzDBxg1Ox2xl7dQ+LME+ZmxWErBnpQ3GBeciZdsyp0AXtwxPabx8Q96
RM5uQo84KEwuoCrbVMbrTwJ2pZcFxX2OYELt1H8WU4w83E3ohfpnDMbtqPs232dk
lVn8cdqbGmZP6ztC46ERBNRA+lKGLF9cX8lu6wROGUzXLCvnxQIZtMJo38TQDK2N
hc6w208VHUcD9a3Yia8gr1S2eC5V5UoLzvfiYqb7FpgqR8oL7A2sBlqTf6ZJI3XB
EW4ZAwWEB3difbKO228DzA7scoFbvv6/4mBlV20+gmkOB91bzqLAsA1aiukdjero
wHJ07Bh2VaLKVAR5H2bKYem+u8YjcXH3L1Ps4s2Rj8TH2UaSLUIMesuH121wS3en
pWcI2GK5P24IQWlXbTwtABbWNa0AIkFjOzoFuSqCNdcLRVw8w4IvqXaaNWP90oua
KCamd2C6+ehXW+kwjQo8LyauN5PVc7UVUDl9bN47Kc3i8AOShuL/BLa7IwDTBWtV
gTZLxKJ6RrpI3t1/ANhkEoQzcAPeB64r0Y1v+vHSrRvCeo1FCrhJLSqPu0RKibWB
jJ3K0Mw+NID/OyQSbTmVcB95Oov0oauVmBjgVAOq3jjxwqKiC9hLnvHsgI457LrK
BjdsDKlhLg77FI4MBIAImXf4C7ff6aZ7+Js2rof8A3lJ6vBmbvSYjpjNxsW5KVQG
VhOgzpzNzpnuX6OUhUq20varj2C1Ne2GFgXSuk/8Zk+l2uMP+AJeJFsHx8Ri/ND9
KAL2W7eF+oRPrAQUJmHyW9jwxWyYttDoOifbxmmhS2scx+iY8ZzOH8+6bbZZy56n
wIGPvVx4miLcdfwB0xhRSU/cQBhm+5Lb3kODeeKEtYaoBtWOZPjc1wtFblge6j/C
DgushjYolZHKvkKPKvcVWjIDNH8poLQS13WyNSzahS4lUG1y/3XJrFiAjetHNxy0
`protect END_PROTECTED
