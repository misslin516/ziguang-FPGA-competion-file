`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HiwzIttg0yFFOt1U/b7TvpYeqj+vRiL6bOZQAuRW5jOHSCQlCjGk+PcpiCZQmiJt
npHgX00fPQt7oB7sj//j7JiSRvWU0a/+7RWIZeUHZs1RVgmKFuC4klfcvg19Hj9X
GUXepa4cYan9Aot9uk5UctU4mVmA+qJ9jpO4l222gHATsmV3aGoaCEK3vmySLD84
9Z0edPeMzM031kQxeRvdA5a5D4CvIfI1RTEw6BOmyh1kR0UN2cySiYX0RMrtg1Qs
TIRZcK796soxp/a4jhX96R2zkHuAivpPQSM35o4Kr0/XRAbySe08qWLCFPqwWzJB
Bee1AO87z1aE1CGmaYLvQAjDTXWXwNVKY6chKRtyfVrWeddwJ8279dK8otItJVwo
SiS87jTJ0pBa9SSFv+BjZdhLU/Lu3kbpPSICwDirSG4RUqNZoAkzO7tAFrQDyz9R
y6x+iKgpmpyW8rFksyokW9z0LutooV0VviWeZpbz7MyPVcurKpk9eXCqNlRVzGGR
ABeQmKA5Xp3+gZO9tIyFmsyGUnBiJJSuRwWqm5YslqiBxFWlNWiCDUDYimGUs1Ys
8FP3CFlw+z4S69MmcBemsVVGz9LSJHBBKBWImIASeMykxv25kTAltNT7nmwS/V6Y
muhv4WWpHMLtpFJt0hF5CrVluwV5iTlZxufMJ1BgUbNRKf198R26KVQNL6/D4LvN
R5rWGrvuEHDsZmjiRrzrseyFIH2LIs/5m9toEk/FjVDfrnXwaZDgOCyuqwi3hFh7
05Z2H9kmkhmR9aLoi/BTU5qEyzRTB0UGFJaWBwnuSY1WSDOGK836uCK34XEsuSX/
2Gtg+p4JaPlAsq0f9Qf+gqpJLfn13gxQnsBZrZXkjeLggNZxRsbH03jxlMogk0aV
WqzmQguye4M8m+yp5hT2jSb2OTKNmn977MJWvo2gFSErERxozSCp8sbF+0AnxO6A
QuMx/tYgNUNhwo9Hi9V3bTC7LUj6F0ILiFDUORC4g1KmcDAYIvRh28gNQhKOQaKz
Gg8vJuf1WtD9ocMA8IKKl9rPNhovjx0JoplAoJVHycMH28Xii0kj6IdS71Gpchn8
+QbWl/m8AL7Q23SNxcxD8Tb37Yug73NnEk0VD9+l1buT+dzoyMqRjyIRrPqZ9w9j
5JdiM6qGWUBjPjtTiEpHfgPJjMpiiI/oWfWakf4FJfBdqlRqfUn5uZ+bl/MGIJaV
5xT0H7XH2lmLuHMoYL0JQkXf+LIVrWe76+rg1nB/yacxk8U1TOiX9L57O19Ool0G
FKQt04Di3q8271BhEGTIUfK0CTCcUdW5cvxp3Pq7t3pOBoVjOxGT3dhq71a7dOVC
G58MZZDxvtzyQ5WASooEaU1SPWc8hrpORPFuWzxD3fjotZs44urNjn+a+TiPUQl+
TstT6/4ADaKsGnAT4WRDE+ooeMf8tM8XDA6j+hsOodboN81sdIjgQ91XjFuc8Tp/
8EQUFe7WpO7N8GNQIiKF39t7g/RQXqr7Qly8MpJJeNyWF4qz81mRl5nCs/qZgUA4
3HnEYMJ+h1DG3xcy4rA5Q0SRX9ZwX4gdKLy1m5ksCjN3AB/Jv4Ayfp9iu4bLFfOh
4wIzPE0CSyOSY0xW9rfiYHGIaX9fr5i6awRZ7nl22ab9qj59BGMg0/mORinOoRIZ
zSzW6Fk6cNt2LnKMcIm5etj9DQAAl/Z36m37Et+DOD8srYskHBwrV8+lPt5wsWbB
A4efHVcBm+p4tsaYxieQQeEWFEdK8C0dGU3lYID/smxoVjNea8dRQH4xbOUaO7/e
bkJttADIIQodtsf/2gyGP8C3UzZaXaV+x7zizuLNF6aT2MW7mtvLVTn3xUPooQPe
wq7LMGXi6BCJrmjJXA7RVrQhuJSLBH+mtMkbN90anY+mJnIz9MnOqyZOpMc+GMuV
xkeAFs5XPOVuxA2sBi1u/Z1hgdRV7OQHAhNeAPcx0pWy457Q38w5qBTD2J5e69d1
5RHZLeBYHDVaIgc2JpHq4dD2PL25edZXx9srOFsVfF9PoTfxnyY3mFPNv259YOOc
x3t4uPTXrIvcdKxFWDTi/9GjLIAAdNLfotRWH/otD4xMZJFrLMkr2/Nbq8LRKjxO
M6HEMAtD/dxQzfKjFXa3CSsmrDpC2wrCERRXk0m25Qs8byTdVWe0xMaFe6Ek3ZhG
SgXXHywnyQTfi90mZybZ6A==
`protect END_PROTECTED
