`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4iKRGMRCOXXbCurmuBpIAfFCJulvRzbyyKnK5m0D9Db2/Upgqhkckn/X9MDrNpPE
8PGHQtvfFFBcfqv5NWURzgtQEFa5lSY4POoAScn6jA3h9rAPObwRCuKtDU2dtHRT
CQFSIIkd4jfc5/pMh49lC8p/iAAcvW6onWqFgAaHzhyVGnm3FPTsrHbeue15J1U3
Gm3JH1+heb3Rk2QdQsLFDtSwVTA6P3XNtoqMdJlIM6UxzKx1UDCVbbm7RHM+fKxB
bUmzhqvbDId/95sQACWjuEe9aBrPw4SLh+QFRmoA+2zJPiPaIRO5vgLH54rvdMxt
NCEpMeynD8//0tePp7mVYEXWhxdJIQ4P9Y1ZEDuOdCnuBmbdOyjfacEtglkdhtw/
+Cd/uA5ppoJvYz4UM5N2e/P5E+qZEl+X9RcOoYkH0Jx9+HSE+HERyC07hNED1qtf
ZTuQuqIs+VxC3VX1IUXZ3X6r2kYcRjizF3xaKHqtBrxeVAWvnkh+KH06BlMivotI
NRlr4W9v1QN4hht46iuT121weUUfT62z/rxGGDoHdzpKTwhrlO78FUcaXEt807p2
qWPkoZZZcUOkq6IEqNOSIj1DS8CGVaMbJFipunAsGGzxW443gsbBHySSfeHnIULl
qs4JQsUCEhXYaPb3ojmlyQBtWqBoeX8Jk+uQoiU+cCPRUSA0pdpoKgDL4DdEoxPj
DnM10X5JbCLmp9UhuYRYa1yDap1mjNMYyAlNeBmU5bfXHdVmzEinqt3CZW/TMK9Z
uQ1fYq1UIdEm7LlYwl+6s5J0gNOkG4t1fshePGixDAYf52TbrAFtUJAOR1cAvqhj
PcUEKSq8DFQpnjTC746MI5kgLFAZQz7fg0MAi5Ky/COYddgAX6VEaWuyYpJNg3xU
kblArfHnjtPCy+Bee0kgRQzWn66l5YCB1xYRUA3sGKwy/tFeG4ZALdZHv79rMOqz
SlzdtBt5tcPQGM0nXPJ5a/nVzpNSTdCN2FV/MiLrgsnIz3IjZrB0i8c/pvnHs/VJ
lTBpl2OrElw46Gk5Pb33EfhDV9j3SRIqYhFyb54yAGcBdf1NF+WgHNlMtNhOW2sB
gOzqVbaR4Gi52DvyMrO3TxLhsCapV6g29IzAZUgStg3ZNp8iXVJoC9/kO8zJDK3A
Q5RDtXIGeltsNBVY9tXao5tLcjPitIPbTEbR2WTx8DpB8pAzMxSNRE/VZHWv8+S1
+98tL++XsGBmKw52mdBSGoNpzJUcc2fAstoisgaMbPevCm1xQJEyAeU140S+cVPR
pKehyjMECQ1jRn8Us5EqJsuullnSMcmNfPLTADswm+H/Q7NABGePKn2GkpWTBnmF
Ly7lHu/Ns0tVPdd8lowoypkcxq6YyOocdnjV3vc4D1Y=
`protect END_PROTECTED
