`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
drHODkLjHB2SdDdS4odlFAQ7Dbuubfrjbs4ycYGy5LJh8zB+l2PNxct2EjrDqCAQ
agSk4f3gJF8waEcS2wIqSpj7MHmTKrKofDejVCaPMje7iora8TBqdvuWMe0EpQIL
lkT+AF2wZDpj3RRgw535uyN+6RvvFfViiH2OZHTEvBzQN+RM57uPXnX2IYSI5dNi
/2yZ9/UGYK08Ix75BBVpzfrQTw83M79+og+iLtyH+Ft694BTdt2uIQMZREopBipT
H8kPjyN19+cypa+xhxQ0z1fc2VzMiZffo7l0d9g6Sp9npTsr2PqmTs0RVXWmRpCK
hKsCDq0S6dxprwazRPKWYu+JeZnexzaWv6Wy9L6e8A1zfwr2FkWs9e5p+TwAMa6P
mYxTmt2n+EP0W/ZArT4JBmw+VoRKN1utcKm++pLt7OYvlNI8fvfJCrOBPZIvaIZn
S47Ab2+USSY+OXNk0c3KNZvjb0MQzVSsnOyHnUm+4+bTVlLI2Fj81hT/NzZ+RFLV
/eQVinCWgU3/3LFw49Q47jK8yrJSpXYv0mZij9jtQOc6pvCgTbryaGfsQakfsZlF
9z5vTDd7oRuEZCoqalkGVbJMzM4HDw6S1ck1ApxjED3WZuB24RYxsmR+QsrmIoUn
LP7TdbseV6tYDNB1bck9QmWTH27vVuAApAOZzDQvAjI89oWFyZo2Siy6ZfYaNggW
ZhtdYxLVNENY72cX6eoF/EsWDvsO/2OrlczzttIxbwj48iP21T9lO0tfTSDrGSNp
yPsIyqoYl9jhr9oVXH9gbrdKDrLwmFeXBpJoIJuqCdqe8zd0XJ4e0ChALrFya8Od
2AoVBeiE3CiBu9MaoMMYwgSoVDGtJ5XS3oGy1oLOvzhrvbxldReCkjHuYl6XqG5G
F2hLSqxFVBEOCZjj5fYNpIZt6I+/V3mzptP8tstsvyQlxmIK8+tdEbTakt2fkmJR
JbePArHQjk8xfcNUGKAZwkNeG9LaP4L1keVgvn3psciQD/62cMtCM43iIbcQtkxN
CvywNwVjvNrv+dcV17oy883cmevwx/FDQPRJRUDlvxW87PrJvmKs7G7JKhpgzlKR
zOLXEyEHLXhg4w3F4O0mkkd7oa7D+LkGyg9M5YbIx6HZbhqil0Rr6TBF6iyl090u
hhMwZ9N8pE2rcAKjKLEPfGeLw07HQ/vtEw5Z5hHvW1irDKNZpH+zKKsy5hm2LjqB
KGX3hYTQFTcwLTUUV9CPDnrzD4w/ZtO6Wq9pIOzc0uUIWt8yHmU6On65fC46H7FP
fMUFvWwdkey2gOJ2pTWDh8ySlp+voBAiujUSbsuPw0hqBRvAnZWWCSVByRQ3W6P+
nnweI241+xGXJDxQBBK6OR0qyJh8LkAThSrsvuzqwWcdrnN0vlVFLobxKx2Jinyk
MdKo3jO8tC+ZQYrb+kx1DODzI5VNkEUkN1pQDZCnDCqWTuAoNtp6gpPc/Vp0/3ee
fD32RkiD6aktN9acRbW1VvQMx+W3wxd9M6RZBXeeE1f2pp9qPUjU6IpeKFOBRAHF
SY0gP9rfAh05qvu4bAR8GQTkAY3yGMkQRTj+x8I9TYkjGsaMsXItbTB5qakROGBw
drtSbVKGSa6GrQ+SmFhEguyBHTD4fUw/ln/07waUjsiT7IqsfJlGjAmmmRlVH2Km
KGAXJLupsQSpKZ1x6M9y7kP9rZWy43YtOKbJ+Ku3JJirE1jN2fWYnX++73znPORP
HEJpEfdGsGvVpCVScpvcDIaaEpIdj/S6Fprw9zExzlNs2YiHAVozWUcixnXbJVzY
zziHYow0A7rEI17LeY8ujnH5Ie5AkwBQfxv8fmiHOJFIUOR0rQpfa0Jklkypsk/x
iCQXTbNAgOYzKffC2Mgci5GDS2mGdD4RHjIXr6D9CwsTPVMy25lk7nDAOnYRhULY
sYyat7vrwwVfDp9GDXmeLmsvEiCPdgTbL23yFOEM6d6hkEw3WIXwP+DWz1VnSCD0
vfyFjrDVjooImBcFI53V9nWmWPTVtnIcON51aUu0Z8ISsg7hfKhju7gIZxbN9cM4
mIEZQmMzKcI1r67pB1pRE9AJo5UqX3/k1m9HY43ajiw6tzr2+HYPz3IYT6oBZbWw
yiOKyhV8YXvaxSaVEfTkRpA9FsfCBPe3VdgxZnrIzdDselnR9vVwt81AjSHMTxo5
/OrBPwdHjq338snvj+2cgL/dESZ7YTIws97URhamEwxrrtEDBiyDWbgf0VN9VH35
cnndsNJiEeG4VIox283BS1//X5AA8KnLFDiP261364Z8SUL0f4P/P7NWY/h5cxdt
czZrGaRp9FxiUkv3S6MsF1sccVZsKER8LUNPJw7MjxT9PxR1FTBAgQfS54pZ3w6t
5+2voCxGrM02zWUQKLXMIBjgPef0XH6X8TiQBcLbchwA0wTcRLrFz7Z4tAhUVodc
W36v2vHvKwqw3s1t7eUk0YlvDFK4LKqy5/CIJPsl98AYTB3/SMnGqTfSutKv4SB4
zmRGwE9lZn24P2r2w8EAjk7o6HgdqpHHMmKLqJXGuBPV9+PIBVJ/CAnkXs1j3IhW
P0tF8kxgKDqB3yL5uyya67bHDVR37YYOpuAZtBITU06ML4NVFOT18YIzZ0ovuVin
pu9w0clujtmwqkQw6t77jZfmE3aFNuFhke/HE7uC+cC95gir36pqttGgE3cC/kYi
+Zprqr27iAj6SNmmDVSTBTpWZUBjxuasUhfQtjKnYAn0tLdxlYyQYPYr8Q78eu/w
GaF/TD2GdlyLKzLXTEKE4EiO3WFy6bs3E4/arUk3bvXEMY9/z0dgK1QNarxOBYu2
cYJ/RwC+7BisJSTUpfQStOtPUb+/It0JDilfHQjATLmNOUUJipgY/MISkY/YiaXw
mRkubCPy56QJu+4fd/0wwT/1rP264btGBLA+vNfCGkGfj1mOlj0ZQmGjrRsfZIWF
44bx33nqDA3oT+yJzHj5OnhSlDEcfXy3EdthPQcnMxQ=
`protect END_PROTECTED
