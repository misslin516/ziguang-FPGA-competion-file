`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+egGAv/nAj8KfF7SkjTACbaqV8MhVCD333MvUbb6BRf3gFRGfocisOmNiF+EYzc8
mFXbbF/9LJ2a2DMbjZV/MIn+QGNNHqF86pOyN7RO1s515fMEQ3XvRjQ4pveAj36+
0H+JeLyT2RVhHkjhrPtntBXRDiQtxWVO9WbEc6dbthU48ePz/SrVTonR3eaOv+bI
lrpv2bG5eI8aenmXSLrhhsSl8qQUp+51UPEEhlttTX0Qo5r2PiCJ9ZDFTJC1s+w1
IhNUo05OHIEpuGMzmajuOC9jgb2RnxtWa3/xhOY9XDT3IKWE3ueSmh/vJs25ewX0
sJYfsexPWK8qa3HVn64ISTMP1WoA10UiZTlgKoZ66eioj3YRRfFqE6HNu8Dj4IvE
bWcAdCCd8M5+GS5AGxUSQjLU6YzT1huXARKeAFXNah+LUFTmuj+iDqGuudxUZ9Hh
QSn3rlxDexInBTtnFLOqyCL9adVvQjeHAxk95wMJHQodKi7cmYOBy+MgnyVF7Fv5
po+r3eYdZhFMpxo+e3qkf5uD2inR+thf4QN3SRGe17k308e/nyzx5Q3HObjvwjIy
oE8w1PBeHCiIZ/oVcEFBdYokgUsKhn6uTFRaecrfitakCqWf7Hp/RKN+qxRwgIl+
SyTwPwuShkLLhI3o0Pgu2poEONGY+WwgiIvVEx1pviKNV5vnqv2vFX7tEo5fN2P7
RCZn/dfBFOjlo8wV/XlYAA1PTORG0pDcUZKENgK36sFybtv46VfP4owgjFpd613z
OkOvzNV7Ou818Qh/zyE1s3abrcwXZumj8UzawWZ3/xoPEvuPlEw+ettIca4CSbQZ
mBco4uognSLx63SD2f3lAKMdFETHbGXS6RzbKOXN/2gQeKmLdIN5YXLdY26HcjX8
jd+oYAMEJ+HVtymyFawH0qIBl/EXMoUUDtgAzuF7ILGUC6BGoLHSgmu+4GyMbqhc
nGj59BomFq9mfJpwok157grdOo8ZI5uzTZPqsXHp6JwTwdtzSX1q/8U0/2aCR1v1
y0ssMxnpOuRaGlVW+U8CTfU00l1vQr8U6+fT+D6XQoYZ7h6XbqyF+9zBEoU+jZvI
ZxH+/LB78AQYZwSA7gehoyaqXmFtzSxbD8WJ/UWaH805GgiVqI4lfdJ65XQ+dM82
C0JrCJ+/UCOzBLuYMKurGojj5mO16wHItPjW9MVt6YZj/WlUw+2ZSikfpF8iKwSn
jtdZ+iU9k/orAD/0RDi/QJKSVsFRnyMrN6pWrJ+7u3X5RQYqPXTGConeAjctSsDB
Gai+2MKtkFlKIVQhqre2fwELMKaXweypzYCxzo2Ya4ifRtLe5HE18Oqn+J9bt8V+
452OnBdKMiy4UEJKZ7jDuM+elLGztt59nfTAPY753zQiiMd/k9qLzLUb1e8CE0tg
NT5FjuIfqnLrMnUtUqYnFkdzKrBq7YqTUP9nwVBVA+JerolsxeYz/JNT3+aMavmv
A365YVUXJo1zUTFBt1erOFROQLKqe8VYSkFNHAuAXBfMiKG1vnJho+OOOPnKxIG3
530e8WB5GJ7YK5jd5JxTH/zIJKy+fKqvqiCcR6hosHYx77wyv/eQKYXIqRvJy5R9
og8b5tpUWfvK7V+rN/K3GFzE12nIPURy3DFALjZy0AbopRRCAjkn+IHl6c5JfrsB
TmF1moSVYxj3hiLlOK2IRldxUPD9GNsR62N+Yc01T6OeXUST8C3XIY6SMFRHQkLP
XZ+p2xLN5yt1NuuVZN1zzryNlnpn6lDIpj7Xxd1444baB/KmCREsCQMm/BzFL3NB
wYgw8qlBozAZSdqtwPr0V9bKYMlM9sJbdHmfQ5ZB2DUC6T3Ef5LGrK2/t3P9DwEg
VuuF+ejUBAvK6xe79/79cX/uQ8Lyu+xGaqE3UEGV9wht32DjFTN3bQpK/1YDyIiu
NjfxuNtNzFEQLWjBfOWbNkgBi26YURd5gzaO9eB4T6fP8K3bsn7NwJwtZLXwZp+j
eUWMO9YDW7L0xUonBgmR7OdDcVfzVc8J376IyxE4lwZUt35tMhqCLawBghu5/b/y
C7byDUfh3J+9Hngb2TIRaQ==
`protect END_PROTECTED
