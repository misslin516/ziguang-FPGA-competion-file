`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8QQsyFtL9Y2JyBLA0p9rI91dyOHrE/4ZS2X2Kv47F4jPiVNdZ1O3Kxs5D/gOQV37
N03g/dDnvJQzUybiuNn2ZL6eoeQfEkWkhO42SVhNfYQL3ZGT9F1Kt94zbJeNqNdp
Zna+dT7xiGk44gpRRfxKpV1TD2G4Zthz9GlQPkAh6TcowK8YX5OmLK8BgoAUjvc2
miUcJ5WRMsSs6tFe1uZq4vH8weDSVu6qE9QeVQF5P9lEOHbECv/X/HYrZ0CFT0hJ
XIFpczhwnl8is0xwHO3KwUj8y13IvnMS22HFQ3dMLEn/l8bjtyQAQvA+mltkWcmG
gQarvS54urVAteUU3DaJwCkdyVHWLcklxF7DzsuLKpOPiLfyHhWmWFLciIDtx6LX
5eS4SagSdCDtb5A20JKSKbSsD6Br6SBmUDqoKwfQvXQRea24JoMKHxkw46AptHoR
yiBf4M4jhTMs6H9B/2X5iPE8taaC+5j93iEPi9CfRaJDrWKhMT5cz4MHh/7CsKov
vM0Oshq7jViNwgGT978ph8cWzt3Pkg/FP9Z46dwIhSUtA0ofaPebTEs/QzpaJnJb
2dFHF4YKRfpBl2G2QvtBG16mexNhPIV8b+mJ2bzJdHxB8OLZxYe1BsSqo8P6Ud7Z
knJm119VCVvJdDvOEjXGU3YCY6nU+LUJtg7PoeosjwSbj+cGIm1nBzMq8Fk/6Fgd
hB40XalrDrlSneS5uuSKKHt8S/Utj5Ty8lp+DW5DGiBoydttRg8C1tDKBV3jMzx6
KePsIUqV6PZtQJBFiMQuvhyP3RslSxcQV4SODtKq+lvmI9X7aZGnLdm47Z68BUno
Yd494MSWvzXtyHOyW58hMPYfQKvCfKfgjpRWPg9XHTxriC6uXoBvsRpPi/4saHPy
u5w6GDIEMdlXH6g1C7g+sNBt7a66wZ8eNwoMDRQBpT7BnnkngWXrQt+E89H9AmoI
Ibooemx9oBpyd/GJCm3Zs9Dc93DF8xa/wnQh4jDaxfb+JdJ0BpwQVqPolLqVQfPF
bxvS9iWlh793Y8uJjVfNPXq1a+9AFs3Fu1cclmZVb5tjW63H/BsiqW9nPfx32HLT
5FLQdL8Vy6KR4zmUhT32MtNaEtKvRDZPyAbN4daBEATM7YbEDQZ8lWrWy+o0tbu8
5BQworNFthImo6ytRB+eINi1+4OyWnyzp1LS3NZy3jUoF9O+A6hhysQeq7l5XMUH
DBY3hqFAV+XV57ijL51VS7EUxuulqct3AC1u28j2oY0n/njfEXhMIDpfufYKTwXz
YIfQ9trCrjzow2lmVgwIkg==
`protect END_PROTECTED
