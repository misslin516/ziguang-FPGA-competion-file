library verilog;
use verilog.vl_types.all;
entity drm_init_param_v_unit is
end drm_init_param_v_unit;
