`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8vyh/IP4dQweh3tAJ1F/OVd9PEbZ+ghV1c9bf4OESwPzO1ftV6LR/EAX56vp+tU
dM23bm0sucBr6hhwufVNDEsXTs4Qyb/m45dpRpdnYfeI+3IYajjS0qUBmaiKRndu
WdrP5GWmmZk1icDDPFSxAOFOIr4/x1iWiHH7BQ4VTxrNOtG+DbrEGA4Z2anrKW/R
uuQ0CQwr5dgONVCh9zEjwTx3TDeksr6MZ8ycUEXd+DZG4dix+Y3Bb4fuS5H5MVWf
nbS9Z6Otw/Ic5Szqfk5IerLxrb+nPdBG1U27GScUctQBvvBSKV7MxHSONt/k1/Zk
DB4ru86uL7nIFINrhBlGwLeOST6av4BFMd4ZXKMZQCojhe8A4Qr4XbgYl9HRH9In
FVucMKy96oBmhHxctzZILGBGGGre05f8o5tEVWT8nT6HEnFHfVUv+UcVK6HYZ8qQ
oHv8azWirlHl/YIJyb7W6cp2y7rxdaaKisPodslxIL+IHyF99W3JxYZ2oO9ymPvu
Xl8mbTSpfhBvxmK4eazXTkM7tDv2sUeh6zQAxifulNgTFSxW1nGbZxg/o76l1EBl
RDFJvGAWrRFnISqp7JBzd40FTowqGak+ZLLxsOGiDH5+Krah/5QG2dCq6+FTG2BM
RALUp15ysjWGzPvytRpEADs4KvUX5H4DQh2Riyh+O1a/iN7ptfl6Xoo1/8Y57zk+
Gjb6x0murD9FZ2gJQPKCZO4QovLPDUZoito1syjRRJ8xkdoJswSx8FwvNUbwcV2j
Dl2t6BmlimgK6I7SvPxEJfvEGJfffpQ3/dxfNxC5e42yAm1O58FOPq3ceLHfnr9A
h5E1uDIYx5/fOXY/oFhCfIC3H3Bh5lW7yB8IC8/C3+jpY0fAtoo48qWWldZLBUK7
tm6BdBbgVIdEBZgbDHmP7OpVYAFYewWohcIFzRXDRYGi9eg9brM31JmGKYlzly9m
AcWvyEkZOzbyFRphaDzFdy2263lRRMUgzCOHR2HstOl23Izr5XmkeJdDjEU6QZwd
qOs3PTRQcOA41o/qR+cZZGQRvyK76dBebjIyZK0+IvkEzxL6eZO5EQOHHnde4Zt2
QwXiCiXLSXVo1bZbWc/4RAOsHO2AskvHGMP7J7H0SENuIONz9G8cGyfWK15Uxrqb
urfdupBTNnSOP0wz5JahwtJBzn3mPCcPqEpICKiz4Ef7/5yWQgYp9m0Xd9bJ+Uw5
bqWEFwyRjIwby5S3TMA9QF+VI+swZWMtcljPFdSY9rfAlGBa6XY/y1bF46TKfwlG
2ugATi9lP6K1w6oQOY96c79+pItam6N5zNfL8aWTGd02IGgwZFeHFTXNK8BX5XNJ
NLqQsFDi0zOexwfpmBy5rCoTzsX0i3Y40niPKqddR2P9wZagnV1Fg1+Ya5HpZXDJ
mZdXrhe9vSe8oo6gcQe/AMHMtanja2OM+WjmlWxwpxKGN/A/w9/27HXqmBmAU3Rx
wWcch4Koyufe5Ayx913eqS2l++zj30VAuJ5yT5TiJ6vhewCLkHtl69YNP5cZ+S2k
eRqNVtDxIuPrFjXYR7hbw6z2phC7ix3rtqzn0DlKnFwS9dd5C9FCl4ysPAkX189z
`protect END_PROTECTED
