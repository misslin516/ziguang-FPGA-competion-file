`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxL5RqcqyTy8PUlbfDKeyflpfJl6eBygiZj55h7VG9ILhYA/Ojd70a+CusByjRpE
UrBtoCwVieZ7ovyCg6fQ+dimsBZf95lgNzwR16QwZGvjeFf21PngpaUPwhX3JJpE
R2Trb90fDbHex1x07aX6KXpw+gltu8L8LNsJjsxFgmmSkJCm0JtkcQ572CcIfEr4
/9DO/xgbTSSOTHX2rpeSwkwvqpxyPJif59kA+H0WfLTdQtDaV4iO1LPPts9RKKbb
ToRb3M7xsTevjdDADDd/H6UXC0+AkucnJkHG4SJZ5hivk7/+UTirh89Hs/X+k8rR
H1k1pe3kE5O2JDUKQCwBUXNpvls/Bnf1w5yPhSuAzoslgZCJ0X1DwBCdI1CwdIQF
QCe9coBgSBLLAlFm5m7K79NZ8x4lWhY54G2gBbfzzNpt73ahQVE9Cai++bV+c9Fy
4sNKKmfVnreuTz6x71gJn0ybMYeE/20sjuBSYYtZKhfdbcFsRAcLHcbzV/dv3MjZ
tJJCnxnj1rfCwZBNg0Sqd5on5R0dnox/GYlRahN9JwPHJSwUSosLnZdlcB3cvEbg
n0wdgyLvcIVVJAOOJXbjTTVCJJ036LQBVIyK2lwgU5hkq+jop6UL80FKWhAuyTvs
6bkHB2tSC9wOw91egCFJGUzJMxqgvfEn0OWl502C3PQWP+WZFLYVt+ERkdZ2noKM
LQ0JNQwwcedmtCW9t9w7WXbtHuDeYs0109oWjXDaHqvNRmOJpgvjvhnyit3GMUWm
Ya5unRm78orK1cVGFxaXGuJHnWSB6+T9JU6rDUK5TRowesACg8D7mPnSzA+lSKCT
5MfO8Hh7k/vTooKbVxWhvTGU7lwAhS4py2NThBzc4S1AkfdL2wzAdEG0kfucMiKh
Bd2g5JJ5hvFFGAqrpLVkNFpnRBkvhavbVqLF4MaYr5TWCtT0/sOXtZstLJtJz7v+
ESzDFX/CVmZxwiGks38br0fFm9FiVn/EG5LVMtcwfa4eRYacSIMpVjVCoP/yEbhW
Jw0dYKR6iUOQjNEnFPYMe4acOzwJvMesEW/iJaWS1/qL16Xpz3A4JJ5aBIS/jzKb
sJ6lxmwpk8Q55jWjEG1qFTC6gxR1b/SjqQ3TCDNiVHFwFKkh8PYS4LejxkzobYp7
8qnmZF0I+kwLEmF9z+PVD5J7dVuvTugzjGwwnuufbGR3p2xCG23DPp/bAQ7YPVHn
uapZpOnapmajYLO5/3Q4k1iRXq0NN1v99yDnTpWzgu1QruA6sMGZQTVN6F5nBNPB
XPMXNo4wGKaVikN1BUXUyBVKWJLFa/hLik6UJHX2g2Cigcq/qbU0FQRZP9T9DqP+
ztD7LrS7oUBNIkKbwVYSFZUKw2PKCxM46DunKaJQsm+WujAUmm12ExfLU0uSaHFz
y7wiYixkRV0JzfjNrP9BzGdZTKRgXcmK4EdcE40Rb+LR9T5MXnD1xEiMz2KjidUV
OD+wbfgXu31+5XLPxZvq1TWqL/CK0dJ0Evx2d3ZnkD1oX4gWNlK7PvrdWwTtzZsh
Q5DnLPbS7Coc6mW/2biTwt8GLglBqs+JaBPlybw86Y86nwaDldUnvzFv8b2J4pmk
aMbB+7LMR9ZOu24tw1PVVq0ex5yPAhTYI6O7pVVkteYQVXOfsi5qNB6BU/pnrHZs
s56yT2JYUP0vR9Oy/9Sk5RsMTcfyiOWqwAKgHNrIscpIxNTD42zSs+9Uvx6pyXD+
9KPNVrP+nUgBJWk7+ODR9bMWq0SKrCcbrVqBXyt8YQ+0RZ1QoZDqdw3195DsF+x5
ga7yR6OFVZB1oF27pRUX71RDxqtERwS3Ee43MuZRVl6lbxYZcDp02pbJb5dz8lwq
dHVbPfAIlhy3yP0BVZph/Npb67SFzSbrb+JMVWmP2MfctHTp5dBA6t6tUlC+76as
JeVzqLjn0aH7K8uzLw539m7XmbR3Wym3rqQOupEZ5ZAfpJJcQvew6ShWJgsM7xKT
Bva7v9P3ReyDyLpjlJxEK6btKwXHak5rydFljyRl3Ubk4c5sL9NMD3UsmJFfK+/Z
blFbanSTNVochGefrZTgz+GBPGnynTFZBmN8sYWA0yFzTXie701ojtLrbTptCQMT
QrfS49ANbiTo32SH6dIj4DA4Aweh6NEfn6vT/bMXOl+QUy6eU3OXyEtDDOqzwthf
eNUbshHvvhyUB/4znrIpDZwebJ1zKmTVYfpXx1ZlhbonrBiZkRR0vnve3YBlQ8qK
LAAVARcVl3Rl2a3Bdv+TKMyN+BWlVle6EglgJmcnssxGQBvjrhwN3xrqmkMLHKaZ
ISBGWIKC5woN4/AASCTB0aoPUy5I4cuWo271mIfjaJAsODWgXxPndbKAH6WI9QeO
EIcuZPnkN5tbUFlxI40xgy9HWX0rg5fcrbmsqOt3eTwGQLLH7n87eWjzweXOf8vA
p052mSPj6PwA8/+YBq07EkhJnSPR3R5OZQlbgPhNgY90yIaDsu4WjB6+MGZqLIz2
MvLrGlmFveSDGsXFU38l8fxDGBdcSwJel6F6bOyk+4aTneBkKKwaV3LyBHTAdn8y
hvmFjvWtNaTHAeBJeYHzJ5d3+lS/e0doJjJUTlCp/ZglFCYDCVORbce91vHrFjl/
vgiuCiDetm1y+yTMy2d40S9k7Imuht/jLSlisQMwcs+uVdlPcHyB9K05+ptNNHLx
Dylc++hOhgzSvaUZFFHoHaePrqGiyzzLWAT+jCJqki5T93+IX0ISqCf0swwra3tK
+ufRxv/+TO1jttH9UzUbA+Z8pjHepQTiVnNMTNm7TadhFQKDxT3S6W4bgph5a8ou
8Snd0ypCLUM2YCtKco5r6GXeWpiooBc+C4PL/HOaG7I=
`protect END_PROTECTED
