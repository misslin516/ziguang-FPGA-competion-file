`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elnGDa064rrH6MObCZN3JBcHjwk3Zfjwe2tDU01pGk6uTYYFFO0RxtsWHBgUM0/6
fV6LXwavg6xF5EpNAaDPUq0Iz03Bm/4YT0Romr5RFcgLWyorjdbcv7Y/LHeccMBc
94ZloImfTzAJqYbKSWo9IYgwdszOMUBVwMybvQ6tbINMVuWmT1jd2vg3fONmJslu
os9R2b7MhwAi2sdnhFHEbAFNXLezqKo2RebTLmoR3LnLQwfpUdE83ZYkHkQtJW5Y
ahYiskbjacpmvVs+ZM0rqJeFIMcsQ3tRWKkUT2HwBNjEWKlPc4zT91Q98I5Cu5tU
tu+J5SojqP3krApaOLOEA3rax9f8Kv5U3Vb39IPK/qIdbX8SlV2pi2C5D4XWchni
udPE2loX8gpNPxn/yLVbApUcWIozBk8Nany1dZUUZ/S1IGvPQi7zgta9DYQLEF9t
MKtBafzraZgOoLDp1alB5QO8cslzan1Bnp/2MxnfJ4QsMK80n6LxdrY816wPHliV
76eL/md6VLJZDMpU4oDo846c/IniXgt59aiAeMx0Xr6xtjXCVC32zVAsFCdLfiRs
ael3av9hT5Cxinq6QTC+XHt3zFYM96wwWFiMEF5CqzqqVbAKTq0k3JHL8Hbp8PJx
UmSkP9pQLnTcxXNI1GM0XVGvQFWtm9Ca1Cc4w5D+bY91TXofdBSs1vD1IYidnYGk
bvJa7fOh10T9Z91rYQGVtdhSSHAnoj+fyCvHadFPeYqT3pS6n5BTiQIifecY8nBn
OavbGSDml3Nlp2vKbK+U8mEZ4M7WAU1LwTesksxzvQ4IKrpPMN6/lP8Ny/QOmBHy
QuP6Djxvy0XkMpHJv07h5fa6LRXN+v6eddFd4IAUaSMdr2j2ijCj6vefoctewPLx
ubtSxTAfn31DKkAejqjc1Hwo7DJHMnnyyvEzI9srOuQqWvsthP6M0ZTBREJZhmc2
4VmZyWB/LLu1ufJ8otvfSHf6tJd+xWrXddQW1dWTY1adZj5lTTxf7MX8e2LQJn3W
9gfDUSy+1c7LcGZUZUxIgw==
`protect END_PROTECTED
