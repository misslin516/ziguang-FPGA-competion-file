library verilog;
use verilog.vl_types.all;
entity ddr_test_top_tb_v_unit is
end ddr_test_top_tb_v_unit;
