`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bu9Cx9cCmTm07iverPqj4rqkB0LiyL2WxieIrLlDxJmFp1h6HPWcPTqeg0g1qLMm
Fb+kDivo7AafmkrrsUFDG37/WPI6CraSmby+hNX85az00guLG/yK5rkN+O/vhUx5
QfoDQuT4cpGTs4ofb//vZxhy/Av5d8uMkR39uVlfzT5UNydyAs+m8swWOgA4Hcs0
g7bM0EGfUGTz+VGaltvKQVWf8mTcLKYRCfNsK3wb/RqSXBkopKN0f9oq0/Q1znnF
2dWpPdcXPUheQaIpNEdIlrMukTqMMU3EFmjB8Xa4PvszbD5S9sANbCc7WkpZvukm
GHf31HoU7OBLGu6VPM9eHo5vH2VfX2DahQbtqfl+60L4i8umb/kYMWKCP2C7pTvv
f33RQZYTB3GUmUOdbUdBLRSs8PRpe7w+byxZqiNyZHYL9I3nuZrbD13iPk62IgeD
Rd4DE9iw4osW6Yi96Dc+szbyeZ19uLlBRVHgjiikPzhUBP8wWhywH/JdRXO2/SAT
QaOKR27u99hcTJIFS0g8dEQmIp4iF2Llo3+7hmsAfi0imaubgmgwnAnxS/vqgT3P
mLAZHhlM01dKV8vNvBXl8hrr5R58cHHB/2b1NMINfxI1oJo/R/+QPo1GljYcGnQ+
g0XMx+JCuc9CpO6fYUB1NA+KM2sE+m+b5vsvYp4sc7xOb4wyiwEO+WRqnFyAHnrb
OinDajXrDN0KYBSHhkpX15Dwe28N6vvGj9aKrVo2zqjTDqjMX3qJAt2gxaQKt7e6
/D2QFogsq7mdqJYJZH9NSmblrR9hrZiX6TyI0fQDoFfkFb92M6HeZQg+zRt5PAEJ
cuZrIIoZ5zmkvn/gzVeywCYgjX+gouYEtSwcjyo03lGl9pdV2V3zV9BrCP/hm4/8
`protect END_PROTECTED
