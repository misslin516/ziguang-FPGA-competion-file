`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1zQsHJOlnpR+BC+m+zi9nIxfRv0t3vY1ITV6hyMspP1w5tZ0k8JhkdwzFHNpIRx
N+xoYc68X1iGZ3Qb0y346ni5LMz52dbxTGsGd2I5sIhXJT2CbG+YB0gNiAU0eBsG
UZNVg3fAE3q/G30vWI4Q8g/cklHap3GmfjMgFIL1TOoqndAVZKgV5j/RWh8U0mcz
HBlORY3YghOEYbLWCQ1o+mvmysnyn45vGh+QyFBMoG1iHY/IpaWesEXVtBGfltxf
jkhk5Nc/+ra57KBJJPAWMEbMQ2eiQHxPiZiUp3liF9/HG8/8TyF1kF2sgaGv6ZfU
Cgq/OeqQe5LSyL1+ju4Vf3JfIl951j29VdpHTZHNF1TrufBmUIdMefipQZHmuKlm
+yhePSDbAcsVpBfls4/hC8xuUrbpcf3NVPm3UKktaSD3qnTlSU3bVp/yHaDMR5jM
QDQ6fj5wPGVJ0fWSW0Y8qovUdfLaFmjYmjI6Z6LXFWxwp7Hsx9J3IAlnjqm7vT90
wtCPznXG1RUyCWK3xQkYNOhRp87QHK1HY4lWvCCxPg/irzLC+j3zmMd52ihJ1Zey
+fL1G08Rk6Nim/RrlcMEWJU/APmIIS1EtdKOrICEZAcKqdqk90jyyiGesHX9i/+5
9fpLT1IvZBrT3SFUTlDAn74sPZ7pDAZJmIa+0zEN5sQz2I2ZeqMVo3zb7D4fkOdz
wCBQ0oHGxS5SZ60DSC55JhDO2AivSIPXeweG2C13KKOffY6n/HMKzZzocFMaa/Ek
3SUkXvEl0pjT16j+3TkPWb5GWOJZeWkNRrX0cA9HZx+QFYcxTL9bbboBndCNRBee
RfyWchzQZIeBGcySgD6kwjMXWYxG+0SJmbOxE57+TCvrWKpgP2QvhpMrfybpuFDd
9dWco3jSrNvtGTCh/u8xGwNXhaYbkUPEOfdZTFzQR6tpSZ293j0IKo5ydfSm8H5n
FwAWnOHmR7QyozOuyKj9V/1roHQiLED+5UJKS4Q0cq6IUikTPqT0Q/JSpGlcAHeg
w9rNfYPoyIhQSfznD+mB+Z+LKPIjyOIs0I4dASZnMxGJILFO+0NW/ay/7QCD0kJH
1VTn0fOK+PdgJVyUsgi1bU07GvBe1dDRzt712+KAINLBcJIArjpmjnw374VzvbFz
JN1+IQyZsGKGlQSmioObQY/gaDc4tRwNi+8rSAAysfvde+AET9W1SBAx4PvAuS30
pSJERcMTc9Y4Vc+KKRFSTnoQLDvelgrTPP/z0na9sMtOrdlrDoBZ+tiWM69k7l9B
+h5/80lfDfAXhhtfflHXtpyrHZoW/StCegaLh6OrGFhJXx9Sp4s9AmRMcvI6AthH
luyAdtycbRuPS0CuGYw7mSr7ypbsxBaa3BV8YAyPclfFg4lYK1U+eJurokikBgeU
CxmbOHrw8KchsJB0m5VhV8ctghMyqDQpFChM4oQowmpoamIHCpAmiRNuwB5+1xJs
+F7GCIzDb53jVfuaWe7iDiGM+VgXwqiv0h/D5Pa3082bER3WhRoJvEeou9KpMbF4
LV+Kud8Ir7As8sdOi/gtQYBNAOJ1QKjjk1B37hlt0AQQE0te50ekxXJgjNQA0/s6
nXy4hbsTJboUwVgC21/7+wzU1N5Oc3tqPvW3DBP3Z0YDnIaXMVXS+/jkt67axKGx
AV7Sj+UGoB04KojZSCck+oQ5zKKCmXlAXE2A0d/WHgI/pnlS6vb0IyWikaViqsmS
DRIid2SK9s+xIEgyRXmZjPcn4jg05Vx26DTal9IwGSoTDSrYx2dc+kmEu2+lYPU/
u2o0luiN9flncrSB/kT1xzDD4pei0Hcjf8Di0ET344kWfMiYHaz8l6awUXaPoeoe
6NjcXe3k/DbVtc4xvXxMAS/9vEyXhRCxT+qwr0pWJzFdkXx1t0rzlUbcMbwNM1gB
PTYyPeZDMt18iQvEtAb3rhwnmSXYIIVlCByt7riQ3o8WnMOuhiSZNXF8RyBosB4g
k0w0sO8O0gGz6UgMl86YDnlBEUgm2jGz6JlxW6UjwEl6Afdy2W2ISF5QGUzwZ2UY
2NndjP29cK/PIRZfXZuTPzO8q8L+qwbbSl2EDhz6aUaoJLJGw2S7To8frCkLlxOU
yTYRAKnCszZslWjaKV270Yb1xLYWUGm37WTaJE4YN0MUJ4ANO74QPQKtHKo2pALy
c/ScJtPqygZ1W1NvaOcDH/Eti9IJBekbqO1qAgNX1pM1SZbzpWhMLII/gfLozcr1
NyZlVj+HarjdT0oaKCOw0KpM+24XiKTTFkaGPYpczsvk5Y6WoqJnbahovKadhCyl
MBMHBUK093KODqS3w3ItkG0ZLH0RnNtftRmqwuyFukYF6ZfLVqWN0VYzYSg6ne4l
nEwxTHA+Alnv6gdNCHHZuhzjsH2Vpy0xSYDKLEv7n4YP2kPVnAWU3deAIZztDDn8
vklnvMMXhC9xUl5qopjaAI65/jIC6wbtLS5IlozB5+LhcaS+9+LJMdGtKVUFn6ny
fSiUFH58XMXz1a9YEJElC4kQTAd665aQhCNdmyWh/7QQ7OPTisaIndZd2JAvNLfz
TAJsYsEoVAX0HrSUaKW+GTp+3IMy8kadcGuW91uBqpvqFfh8376fFccK9s4Bcung
Spzn3RozMR4E3BOUqvnEEYQIrZ68Z2HI1Mw3S/lI46sDYu0nFV64ts4fEjiMMI9x
P2nzUoyPSGhmC7V4OTc4RP3UDoyE9cflt8twibORdcOlTNPH6BMK1kCCmq2p+J7k
jYcpiMjzZWKZlnhPWAX5yWj/rWXsJ0keNd21VqOaxEscPt8XuCDajDFNSIHrtmBK
w4I3NPmEsv6dsrlW0uJezlwPH+4sK+MbuxzOKrK8tNcwJ3s/macJNIySxQB356f2
/PKISRe53F7aFUbVe78XXA==
`protect END_PROTECTED
