`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRm7A7RN2jMs67YCzIeZZrssiaU9b0QbdDYlgZjyMJNrLxZj29bZ8+rFD6UqxU9W
taSYrCXjIp5wevrChRvrn1d1+v8kWwAOUAeq3COYvHjDaUOuRdb7mvfgbUSQ9EA+
k/iKYXW6k4MSWqLBlR70cCbeXcWAaHjH9BodbckG3DN4v9tw3awPtlyGfvfnE1wL
qpmXuQCNauDbQG/v8REiLItAAsE/pFU9IPFWFIG4hsNTHWiNJD/B7r3yZhBD4dhP
xFhRfhPmzVUKB2bBN0erRygARoPBolSOqCWwoyWtPqUXHuKtqQqT1EAfhm0uXFVg
N6zdyrK/BMK+nbuYen2jQYYWBzZYzj3N/osw3jYXzj2qm4mtxadA3Tu2YQRsYDP/
mcHhPOJJ6YSrMX2CIVaqx6BWMGp/yBONXTRRCBNQAMJ2AaCPOj2bsiOZ6ffoHq3v
2WkA0/4mMYEeJUChlVF/90miIlJoV2hLdvhrcnFl9NLXvYT9LcBeiZb44svus9hM
DTpytMw31fv9uudK721BDbZ7CWTHouQRuLVZQuA0bERVfsHFAU+KskJO7djFTGTb
3y15IdA6ApVo/qECNam84KU5hzFOb8VFg8N5RATG+r9HmLNFofB/pasPtKyickAG
ZDqTYV3UHuFaBWPS675uyGtQ3FvIwx4vV10scfCC0GNsQm8RlqJ2fm+zKtM7QAvb
TJoatvOyahAjyj2PdL3TqaJ+sTBmwiCMTfPS/VL3FeKYM6jXvSwDSYVsCdqQ0Sph
sPXrb094+22YyGryOYh5QnEeZOfowk8B5sY005lpWCY=
`protect END_PROTECTED
