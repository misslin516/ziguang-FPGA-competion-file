`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zoijGyEf5NXGnCLGwzIWrPJgnqQxJiiUU/284sXACDzfYSGyUnjDO0ylVk7i6tW/
fFbsDYQuNXbt8z/01QJn5CvgQUqrLEmfWXBsRM7gXcyW5dfnKLWTq70occl5nY7h
K6cYC+8iWjmj+vWc7d7mHL/5fzPt/uVk92RtrnZkWhWzJGZPS+/DFiJf4DkhkoQz
q1R4jo9S6cW+QUigpIX9QQaytIQv/H58d7tvGFVY1N5K2Qi/GqJwH8EoqPb09kDf
fyoKr+npNjok7xCyUyQ0BEkRFAabc23wvlQd/+4H9Re7wU7zmPo4tubuS56xhEsH
CrsulDvYc4/9qvmM5N72ClHh1V7MmRzpgJCWiOs9+S9Zaw/98wTeZx4V5o98Wai2
nd4NLQ9XsHUhRnCeKYEAvwdlgaC50WtxD7BIreMxjjthSmu+QrZJC5vw9SCcnXal
qxOdCp3Hnjh2MKe+kumLobs//IRosGPWKrd9PLiONBqnUwUdrEqN9T9BoEXly63n
ead+1BEaNLsm62qAtrudDOzjZ5DmwhkXqtvV8rY4wk1tNRax1VsLF9DAOnEE+3GM
wKp6H64OVw3OfBZV69LyT6pQjZUlBLCTe/usEaVwbAXuBvtMdG++lucgoaLZhTb8
kEGKDE5yjuMrrzmw4Maa6CNXRBCzxfdJ41x/y5/GB254O00AjQ8SQ0yqQMfonPxs
mQ+mXjnzXq6OGJl4QpOr3Z8dQ7JA2yLAoEftlfcQQMiDxRb0U5QBM8sVkhoH7Yvv
Vm5g1TcuqDawdwmYN6SiYxTwEz6kk3Eaht1S2TpkR0gf2D36bIgtOtG89AXyGpII
s3Mdmn4R6WcLiEKixPtibcmC/8ZIX9akhVc/Y3GtloSF4yQHt5jwP5/37Jcdf6sk
F1ecvS6fLgP41HRJqFVHMQR+yBY+HSxOKW8jEgys5A7TpTErnEDmN6zOyE3fjNB8
+FvkFA+5oXXE3USQVtWhrvw//ICNAutaSMYzGmzbqXdL3OZKwr2Rqg+DvAZfB0YF
GVYX2pqoJ9HPCDtQrhC6TA==
`protect END_PROTECTED
