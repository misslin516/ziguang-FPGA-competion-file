`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TqkKsSlCJ47ljnrZDP2BV0sAUE+vREBfmVw6Y05RvvZ6YCtCHHCplREykFcmsEmF
Wnc8c22a8ZoS1NLy53zkM2AqmgqjD8BtDEdYfzrQD0jOH7zKEoRKn44mlmeChb+m
hsIMF8zAV4oujghfRyN0TvMVJr9s5iWzXP5TFtvZkQnQ2RNtSt3r54ixk+kKiIjP
7IQBVo0bXOsNEJFslhzTL3YiP4Bm0dAYro40ox3wpomG0n4IsnvixyKtjyFqh6r8
nFxbz5nDLPGrnjOjqugEt8R9UD1bTKtmMNd3ZNhEY/EI7xLY7M/hFCgkaQHD+d79
srSzwlM4xX2GBdzvcb7u9mBNs4rmjKtQBcJJRCMHQzAWjnHDrBHDXONVjbkQgiJ/
49OcY3uWJOwdNw6Zy6qYxvzauujN6d03Y3CgFPZanntSKxpDkFSb57HLfd5Segwe
xzKEozQLnSvXeEL4S0ANyyxyubFTgABnwKl17aXubB+gJUXH50NX/0unOvoSS8gy
m+xIB2+8MFN0Dg8h7K/MIVbl6fp8rqQ4YxrI2JUtVGo1FYSFbOBoEXwzbfGb4yBs
5AVTIstlN/GCy5bOB/WeIH64tmaeeJKKoGlwHdUn7712dHrt09ctZ8KzIpsyEb+p
fqLmmCA0l2d/U7M1iLSvhZCjcCNCkihLbHQgHp+fa/CGucaAO7lrC6tmatOsn1I6
+ZyVSG22kSLs+SsymR3/41asF7WKtqQfhuFqODyNYYIC6AskzuTNwjWCIQBEZrfo
nS5cPn9knXrGugJ5qKeEwpG/uZ5v0ywprtMZx1GnxojsW37yvtJcD9bAdLPmJUC+
bajMHbNGV7LzPwerLXO86K3155G2qNcfz0tHJqpf56mORqUolexzaI44apRSWnox
+2/4cEMP1lxydKIKwObUyqGjEnOyAaDLhFmGLk6ag1ikSBGcshn64lXvs/hzq8MC
pRpRrElX4v3lyIeLzgPyz8to4aNKBBNBGPnGGWzCuW/67TL6unD1AaZ26UQ6eW2+
dc6zWAoLpYqIq08Rsxn8XQQkaJtad9bwfly0U1VhpzgIBTqAMPhsCGJWD4/Ihpzd
j6jr1IwMxmtJsrYQaClY6ZXUZx1yIg+SeirhPoVSXhoivFTe3pIfmeJ5abhibPJ5
x+3F2iCnc89hqtPq5Zh9Zi7BsqYuVpdPXnNAdvuzeUwevSL4B1CDk9r3yo/Pwc4w
rWMoT8zozK7CX/g5Grj+IpeQ7UI90Iq5KDEXyN5GLFjf+ANdLAxXilbUnjBUpSCE
FFGPEo1ExTf6frMSpivVw3bjHRx0MYlKf4KXHIg0ywc7fy0Hi49zkfnJM7E3khOW
p0jf6let1BM3s7q+VAB0r4QlqLsrIZQWVAQ4nCoXeQHK/56YjjjVz1jFaWXhk9Iw
FK6QA+0EESsv3GFQehiV+2AHjoe+BDtcYPoYB/e5YQCdq6Il7wX83dzpPQPiyqU+
8vF1H6OZwGE4JnTc7W4MOc8PZZf9c3cHX1X0o8NNx/oKHdjjf9xIvnLDytXI6ZA6
T5GG9fpKs4tbnuiiHQsjkKK2qo05lvpPCD5TcSMLZ4b/DkwgYslhkNLM62E0fvkI
UdghAYTooRizPAs/6J6OeLnE8Roao1Bda92VSlwKEwvyQDEfbmelQqobVrtvh8Mb
+VbKjDEvzJiiMcBamI0nRfaEVcMJDPCOWv+kRNobxTMGlI/alfnwQreP9zqdrWHO
kOzchR2aVTmkL5xZ3irUpOFy+CBnad7x19lz00iwYF65wJWtcYgpwPDbpwAAa7pA
h9XmAKJJEnq2gFZIrppn8dObAXyt26bkrO1mwH0y7+RkDqWB1X0ks46NXCbIm86s
vsRTPiAbq6PnMPgbYVII46VoNYldRo9MUI415ykYtxPfiKq1iV4/skbRejPjRDty
boJ2MHbZ6y0yLYTufvfxsRHJeZx39jcXoJ4a83m841EUif7dwkM3NBbjXdtoZo9H
8Bai0iLYQNwQ9Nfj9xeu9Stu0zkjIoWp6Z5jNFJzarCb9EDWOXjlLukzjA7p2nYS
QrWHwxivxAzhubURTrXIUnJvuU2t61tB6UBhcrBn1+ekJeGV5lp5JMvu3c5HUUuC
PH89qLWVVWzf7WOw5stm5oY9Crplbt24WhSsUCAvLl7SeIyyYmW4epCzB1wz927j
sZ3qm+7vIzTm/Q7I4+VXGjTGOtFqbGTQX9BekrljCYdfcNExehF3UBkY2Z0VjB/6
JYxyf94oH+VqHZpJizZbzOoJMNOKbINsc7jjrguP3GdjHunHL/zf22GUZFvI6ELp
CQ4PlFovyTX8qA7s0iTpOKspoF0/IjCAOrKceUkHOe0ZOsdk6C7sIn77gRPkJErG
flrc7mH7/yUGed2DP5IblhkLLa8xOeqkhgYgUqhBOwFiol0ElNYB565VUkjwCLQG
Lft0HPzU+m+hm7U02uiR/ubnX8ACdR64utZJR0lnz7O37qLyzC21mix+aH9/xqMq
sJLJwzRB7x9G7aFLCW10BKcgweekM5mrr0J1sAdem98Uv4fCXYLdkCBabFgsy81s
Gt0QPrWO3Nt6jLBMui7moqOvX0ic65g+dc0wkQdNFiW8UKgRODMwObsXV9dSdi2w
Pg6+njgydbGoeKkOSgYkcCaysdgdsZHQ2MZHrd5kY5hjs/fbNOz2VOC2zvBQSDre
kxYtHzRgjIrvopBjjXz4106hBeLi9DBD7Ru+fVWRM6eGSlDUczAdJIXJlZcMDwEm
GgnPUu6uY44xfG6rNvMBENwI3t3tR3B+d7bECpGHEFDyOUZ+x5F6uHXY1iwE71b6
2b2wsAuUVfyhDqCTX0M3zylf+omRFFNQVMy+jR0jL7s0h0mMi+2IIWy8xgpOeXlE
lsI5XuvTQ8jZp801EdLcNRO7hZMvrz32BekfeF2/RgU3pp/FzNNQyH4npeF2mnKP
v/nPVU4GGxiaejwjHl482MMYUGfRQjJ9RPq9BZMYoclABj13+U+qfsW/AXqZGJhi
uM2V3qNJfDSCSWrcAq2o+TCWdEDgHjggS4xZWtKBFGmVZrw4M1BK/pulrdFt39pV
wFjVBV6qYM6fQs7LouwqpmGO9sOwN3K1G8wEJDTZ0wnWh/DQvHWPaPXN3s3gNmxJ
D0PKextASPq/sTMDSakRtR/zw1wZcDOJhS39j/j9ia+iUq0yOWPZEpFu0aQ/+F6a
uWj6BuT0LjKlsRSh0aA9//5LaqVyTp2YCszl4pv6zCXgLIB7xRIGoIPqCadAq9tJ
R0MsZjVHE7GeFczQuf7wxHBaCGGw9cwzua35O3Dg657YWfxATCOL1hd+p4FURw5T
9cqpxbooIJzSdNdKyUm2UsvFrlcKvWX74tnCzi72Yss3Xz0buPCJmjYxnwqf/DyC
u0ORUwDZNzREmKdQ4jKQV3Au3wfzZ1MB89d9MsDPYNKYKDbvQ+h90vR/lFOUllPf
D17wrSq5Tjkx5FpBbAS09r/S49UMQB/1HrELZ7Vq7AXI8EB2qw6r22sXo1CZVzPj
My5YrCfaSXx7c73xfOKvMW/+IIZbHlQebF0wayr0li2+MsYqXxRizEscQRgequMM
dHc2E4tv3vtAxAFjdKMzUQQOdgDCgYqpX1XdcBpe7fZ0pHJbqAz3iSbVCXVWcLff
KOBOV+89Ez8scCPLcmOCtiC0lIlEBeLGjrrIPI17ai0=
`protect END_PROTECTED
