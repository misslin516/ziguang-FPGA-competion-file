`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44tmDFKhN+abf39H6DJcp8OUeNbFLGSg0ii2Scjd0KBnDIw+287/uYKDdtIM8gBw
AVEjLWhvFO5u4Z1luCYGLzDm9eyy52mkRzXOzPAm8PL6hnwn+oyncTudHTt6gILr
V9C2Pj3rBOWOtIisU1j2DXM+tVms+U/3UbDOPmgWz5d6YJswVBw+iPu+qR2zEqpf
NZqqvnUpHX5pVpf0ng/3pbmOZm/tCACpxuLXp/zNTi/akGJf8d+j6YWW+DxKHe6Q
q2DouztJeNi9gH2RgLmr0hJwnU7TC91ELOU9Wc9aeKjc5YhB4WPtEJ994ZtQPVEk
Ne0PJ54iQ8Xcpka7LYDDPE6486nMcWpHNeAsfyduIDWBeNPK3Of//RpjkX4B6bN5
8/3IA57v3tQ46KYOOf+MUpPqAI0TxyycIE2SMNH7N0BfuPCUC5tEMWsyYyvjB761
9VaL4ksRhtBjYK+9OF3XQ6m4ZNyLTTPqm/HkmU2UlxwVLQMz6bC3WcfZbbfPi4rt
KAoV4GjIaR3HDJH3ex1I8dLbPTT+MR+hXlqSnga9fUKb+FxP5Tw8t6CHz8ZysUJe
lFK+C0EHc+GdGd2KbB33z1p9SeXJD38BzYDaAOR7ZH49AP/qTlmh+bxc4trkWnHi
oFiQQ/kQ1WOEhU33NJzaybFZUpDgN+Ta8Q4vEVsMMhwu1+E3BwLNVRI+9dCfTGuu
aKNasEabdAY+ut9pG2Lb/7OKgEPrODSjQundyWGR8sN6vf+OP4v9XhHoNXq5qkAs
ccgPh5b4IXRPl0giiKTXZnNXVMMy/B2bbFZ27uxHpBLE+MW/Cn3icTRw5lqbX4X0
aiuflK+C1OD9q4waLnA9kaXGx5bJhc/27mrkwVuyblAOp5pjcoXOq2qbdreFrLte
u7rnJ5l627v4Jt5/2w6vYvT9m2BDUHMRnS1OODZ3uRj5sys+nKWXUHtPU/cyg6e5
vj0XurRkm2tsLRTp1QZtkNxbV1aNfEGutUjc+em48axT190UJPQxBsFIc/tllT57
iqRUJHxU5hAX3DcZp+llbQ==
`protect END_PROTECTED
