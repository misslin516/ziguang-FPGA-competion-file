`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6uN7q3UkNR3xFf/dltOpQ/KAAcyYJYu8KqDWb8IaWWboW0JPW50YU24um4e8Ta7
tTg5ihEU3NbXNU79LK4KTZ3mYFZtvkKtV1UThlPpvLDKVqGZ3yUOMtDNukGj3u3F
VEkPAMuLUhtIPTCjGFU3ASLICh71cgpVkPqq8m3JdJptO1QCewvOm27OcxiXwYkY
rHLo2z6m3Xf7UEYhSFijiHy6vEk/dw0Fv8Kp/O3rQzXKY4FHZxMP4Krt6jmNXbXK
57zm+EeGusdH/CXRoQg2GSSuzadfZhqqAyhyvaUw+A+4TEh9H4QRd9F+lYWuZ6zQ
YJWmFIqvvXmqT3/5dA7mQxd8J8una/oUGCC1WsNLBkIlelVZNNJ1TZoB70miGtng
F+gm6xF0YD+5nypjetbMNkb8TvFnCVP7aTw/n70tOw4HrjZCrmadyKBftTzLO6l+
Cjz6ukptWf5s/q3ouYIt7Y1vY2TeLIcxkla39IpzAJm50161LUFzYjpf8jCFMDMr
uAPOs1RuIGpQiAh03o3KzoO4QW2krXMbLsil731O/EosG5BusG8sU6Rl+IsAZGxV
xUO6+d6LChqVqv/B75b0IPq6SIlk7EWQoXqkF/e5Ze4bJdj8PMYa1AxJcHSYyHmx
J+PuM6bfWKUg6hQ4cPnB158pKGdlEiLOJrjrwBq7wqnYXX9tFq7p2/LamwzhCBcU
A/X3UliWSP4zKX3f4uvXokg/ocvGQX22X1CjM52KSalGicMmZpUIWTH6+RbH2WBW
9vKAVpGccTb1vRJA8xd6eUblScFxx6veAwnVCB4ydIeUQ0mE4H0BsayJZhcm11vF
5qmSdo1pIz7ibpUoCmtoLKF/d/nOA8Y+zrsF74BSdrDcfcSatZxJdMvadit6I7eL
DD8nMNznH6R3gaFztHv7OrJDZQJvUlkMC8uHRez+ToZrdV0s6LGu1Bs8LIVjKvvn
HKSxrqlBNPrIea5j+IGU9Q1ueGU8txPZONd8F/y4YAzrYFfnBCjLCpmaPgdlsrvr
PY7MiuhSzvT0i2NwR8PmVfyPnbpVpJHjeIT0/h/+4OEvxjVHdBHw6BP7NEVJh3tP
siOt2Mh2fiPRcUlTdFkNOXuzxTzAAwu79zlMFDVDwXyi6IcSmNw6T8vA0B1EpPAA
JONQ3VDYkLz+2chMD3Lqf/15/NBoNlec9FFs1sZh6X117n9VwhobqWW8wYOCxMQp
aCC7+VAibAk2vuGj/9FNb2T3vD2Isu6RMfs0q/6cKBHbjvEY3m4hynYSwPtpOx0n
Rv2L+CrR65L4YiI7JEgdnnsXCKIzePWuJufVdxYNL7Arh+XX9qFgAaWjqUrJEh4W
IY84FhLCaEQqGQHmVlR9NTLZsXhhbIaWHAQbulxyuAhwWIJ+VhDF2sEP+KGWg4iF
o3otZWzJp+kdRFs1xKIY0AaWkkEKmWX6Z3stJiNagH9x6qCUcoj4eMqU3FKF+B5r
Va5fKOlGjE61lsA6qjwTJmbL393Qw/ujqgEJa4QiZUXja8DkCSAaB87dFEsiing2
TzAN7ZvaFbtnwxM4zJIGNekNeFLzchoMELq4j7LprteHRnQFDMoGvG5BLTDyDzhd
tfKY3EtL+CDpn2ETJozKdRs4uhep9cAMVBYq0JXhVq4omjm/J/J5j6pGlXDARvXU
wh9VjPaIbDlAMIPm0RVKNLkLX7BZiuKrml3OoOrrEVN4vzOGCe3HU2ZLWaeY8TUO
oIhE2wLdY8p1y0iMyFoIyQudOzyrGMfg9PPPXt+Q42aiw0dx5uq2SW4P/rg01C2J
tLVpC0sMP1MN1JouATiRNDQ0dzBG16Ov98xB69NJvNKi0jn2d/QEoc4xh09qGVV1
VWfI7zNZJNQPfPcha5PPLgS/M5mwYTAKX2FcSRkIZKDfukuFTGCVhmCOnDCz72qt
S2K9nC4QfbypwoSzquQw6H/a/aPYdS5UoeHH/zFcFFrXjq0rMAxeaHAeAeY3400n
HMT9gEERGFssTLonEPeKnUA2U5OUOdiHLVtplVO71KOM15MSj9fpUpypCX/HYTan
AXKohV5HUE4uN3/wTEGHNZiK0PWVHFD4u8UIqS+JnIMjcAkA1ZBePaJ3vDW/BcEz
EBt4g2QSbBjCV9/HAV24894YI249lhS8ruBo6AI8bllqKgyJXPx8QZSel8rCAiW0
8tDBMAlw1oj5GtyyETu4+XXvyisNJmu5znj7iwsjvOnN/op1orztwsQzIzBKe7YD
QgRtzCZyNKPTXhypSCnugCCOis/JgiE7B4XCNx1VWSrQCbEwWqSQSEZQ66l2bNex
ukea8Rb9RwM0fiL93E7GhjucKBlOpl2zZciyJ0WW4kULK4l8D2GQoXf1sn0hIEv4
qtVNXxMMJEbPUUrhdn//XtuT/LH/zGCFb97KwAGTpK1yv4erPU8v4VppIZYG7Lgz
58GIDNxDyOwAjGKpaexDtcho3wB5gxfdU47Ks0IQbSe3tK1FriB3I09udpGPXR5W
XPXp6nlqkHGUgLHz32o8LMk2vJw+N6iklOnE4Oi80mip9v4xkAab2id1b5kWC8MZ
D+BNcPq9MZOOutVxQaNfxXoSJXFYvVGfR9Pe/NI7RhPxIx2888sdHwr8354kA5R4
bC5cwRUOPLWKau63IHTzwm5YNRHJlgIBk3d7S5l3MvcQXZWAxBN0dIJh1/agAcaG
shEmw6OJen1p97gc0UR8tlM4s9o4rVYqSWrq2UbkJOirkYs9o96DZhk8dw4hAWR/
imlb8gNpeHxZhCo0UO4pd5xmBQxEONRFFZzCpY9q52j01eWTYuYq6AX2ZkwHpO1A
DbhQXvIeJtn8xCOSle3bN1qHaN3O5Sw9HeiwtnSFN/wBxnz/6EGQo+kfJq9AoHNo
7JUcIB8Ur0x0/0BDC1IxWFEFavVyD0ycJSzyX91PLiY1Kdb5yzoYsNY35+roRy9+
O8xGEiAtl4vnNIVnO8Sz3ddHElxYJhA1+wTlZlIJGsbzpt6LrikgIt/FT9eb+X3r
QD6sLe+N9v2A6+sD95O1jMpGo2D2PCHYGqJi7Ot6fRAdeJd41kYfgvR34MmHodoU
xvEYe4olCqL3lpHXNYEMtGs1/eyULlP8CiBnAxLyFCLIn8mcyXWaVk3DjEHZFwsL
DzFz0ajZ1/I+FXe8NUSuWosRWVRjUK/M55nQThjtSeDG46Uj1ul2zL0xDipRAG6n
dC/SbfBWMYHdvcTG2ByvPvJfz329thARAgKoc64Xce9z4IJZ5biPfhTf6RO9lu9b
B4/vcVktHAgo5elJ9xV3/f4KfQ27zHla1bD9OyONYgKKIs22PL8DxD+H3aX6yhh9
Tsl0zoFGlao+hqAe86FQZl4ih8ZRzEhPD2McHg4lWRxxVWH3WJTOpAz7wR/VHNgV
DR3UK5UfnzlwKEdjY44zxIaNKuQHhZ92Ze2q4Rn+VvP4BICMcMoMJ06Yy7Lj0hSO
G4vfmppl4l9vV7TwqQjb7lBEq7C3+V0F8TjvGu83xzm8gMRENMMDtzERM0nsdQbI
p1hbG0glrE0PRcF9jFICV0SEi0OtsbrkPpyOsxUp37O9kwhMDSsapMD47af1Lrkm
dhq50uhFmYEYps+FT5GnV/0kcXCZR2YJpJ/IVHPGt7+1BiFN2JwGH9ZAe0fRFAJB
/2zYmxTL/wjGSvnRmm7i/H0XlVrKb5jwRIrILqpaUOUuzfbLvBfkIjgFCxv0dzqq
EClH2ehcYgIEilMYKoS+7VFY6OrdLmNbJcspZZy2lQbjinuCEICRHulbc/O6q3eg
2DmhyKJRzhEOuoGdtTB1iqqKvAqjUredwklREOxlmLHB+/FNWwOoJ88M99x5ysVL
ba/EkC64POKmiCQzOhxFFNb03sMktRrlGsKuDTXPDeBBhXIVBSqMJeo4h41RXldW
gkcbeVNQkgc53rokwbsjF1lATiagp6qzNsb6XXY8Woyaf6ag7iBS83g2+Pz7u3ox
5fX1aCCJBiQNX0GZsispJS51HzsvIo7lPkqi00u2zm85b0PGFbrl2PV6g85sCWUO
7IWTmmdvzDG0FTz55AE5K6UPfCL3Kxm2VD/FGsHwt0XoqeUjNdV0fbLJeJxuQxow
0rk6Ubre7QF4JLSU3CPRsGN2eTnpHeifqAw2ttpTrEYnNZZSF+JTq/vpbYN0yGK5
XMqeVVD0Ql/AdIV5taD8lnJSAlY1temBc9RQPh2pyIJA4ySiXlLsyyBbmvJ35nl4
6c8UTSxnf2K9HyzwPZOrhxGGPfoH1o21fgh1+yAXYg981hC7OS5O02IPCmlzWkrr
VXb01Im5emOFr/V1aKlqfsqSBSShZcj7v3IAdhlvHhFrBikNQOl/pIvVllhWc+yL
A9sDgr5JvemYFmnNV1zF9Cwk5KaFcjvwg2ufSPIVJitNnVmntcFpYy9zQaX+3O1o
3nX10MNjuFwa0JVuUZCoD0QTelc4/+aRIIpHbUzfi5UqZhY0KYgjIPi02iQUXUkO
1l+2q870r95aGnN9hC123Rv4NlEIE8saC+U6msTZt/JbG2LMCLtp4tk9AcHjP5nJ
XMZLKGiffpXwqvoB50bZRRSGmvVgu/HFvNs47fuxGjk5fbeJdBChm/XGQ8RZXel3
I4q23dB2uMvbCfRM5QsRRisRqyxNG9g7n0w7amrU4LVq7kbMCCnAZ1g2muKlcmag
SeuQSx9LGbScBY8XxxuAyY6qzFmeAJm2s4RGfb9JHXGi9yW7dtG4we2p6Frme0x3
XedtimplZlnGod7pXnArlmvEcfG9BE36cASoUjrA0zJDl+Z1lUOTO1Rr3J+LI9Vz
4JJ6GabVI3lfUM3hkdX0zcczHtO9YxhfwzNmKiz8ddLmjiHcOEoxUtf3dSRKemvd
W05n/bWCInfGBy9OhKhkWztZg8v6LDB8SwUEPA4WHArax+mAUKjB5eQvmVHjnjHj
TjE7kF1z41FfPQEeN4foHwKo4Vqx7WDh/P6ArAYK6GH1odw1bekSq1qos8TCCqjf
2KQCtoBiWEE2h9YW58yVSHOWMs3jsWprInlyVcjVFZwtrbkHPEMAFFt8PA3ixYbc
fge6vnvi/fv6leHiUqH4onq0TeOrxZymQt1+ny8dCoxzZvFa3k24PLgwCdmu/ywe
Yw33LEmI8ANv28ZwtgWtaAdx4bU7TP67OTEZz2c4sRAConrxkBpHqmfSPUP7zzHY
Lu/7Af7aV0VITGp5OXLTqhtNIGzqUQUUFKLgBomSH0BktkLE4hB33zWEjWHWUJuR
wvGcFfV5fEWhDYNJwWLXXgAU8uoxY0zFu9pipZAwDPjc2u39AQZRlCc7Ok55Dq9u
lb1bqGFXggDWbpYxOsVWD8gpY0cJ1d3Dt+L1hAssyCWm9NvQYpd8XjWEZI5D+APJ
fzHPt0jlD/rCtcZUgmI5Jlq0c7/ohzGLxJ9aQXFOzjGdWSMGoHpCoA7v2Wux0fKQ
HS0QBPOw4lu0iheOrXUm6XVDjqCyXvWr8xYHTI5tJ8a7W3ThePTzr3CkHuW29LxR
J/9nFF1ShSrcn7K6L1qVDIAxoUElpqFXUYUF07NWAbXnXYT7PkcCdjAhti6bP66q
ZQxhQhEO2vtTxggQOe0oj10e1hFbwWYQj+eeql1SLXFxzCc7XNGOMO0kS8+YNce5
qZclS8Y5Z7HF8QxIzS4Qa9p8mcf2Lht3h/IsAlE/FJ0l25aoJfLtLmdzlEqddpAl
94xeHB/k1GJTwQXg5tBJ+3IQt/IUKy/oeaLdD3JYjG7Zjg5dJdZ9zbU3DWrG8oJ/
VGN4R4SEFra5Mj9VfCAM5QHI75vjbJ0KTf3q/1v0yEvrqZo8qCUPs3sZTzjZ01y3
xDbL1F+TWoUpgLpWn+gaL2vaRX1MInZD1v8LzBj/rDQ4JFIbdGhcz+U0c1DVD9mT
8hS/8OEbf8URXEbHKNVYFA==
`protect END_PROTECTED
