`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5qhNlfC4W+Paa+S5sDC8fnV/ESINOL2UfiW26uVBgVUZG5wOw6FmY8NquVkx0oJ
fC58qlaTmvOSRX5KgHvV7odE8WdJg/oYUzLlG5r9i9KISx8jAfwZ/5l9PC1V/ihH
QdoiOeK549E5YKaDwihoUwQ1M8jb4+le+YCTy5QDORudRFMR//TKQARExpXVeYEc
abhfoI2OG41mY6kJB/Bd5yawdHapM1gne23H8AgocYscwj2eKTBFEbSewSXa14rx
SUOga748AeJ6a5ooYGAWC4GjDiucWpVOH4GiexLAdCpzv3KGu5SxjyetT0JhuAVd
ID4XlxY9+K/9zJ99G8XO3ybzOqMbN0SSFezRuxnorGdDwhkVs5ttIzYAQwIdLaYN
Iq1ZLpE14e45QGsBaZ9Ih9x1z1XOZ+uZ2Yy1rks6jOLVjXemEJ4PvB35xKR7Ijh+
Hp4Ff2DSNJRup/UC2PzysnZmKDDFoSFQ3m4emLnpypPk/uUOboxKTLpQO8EFzPic
F8WOC3Sb+D5Dq9Vc5d0CxcAzHE7rl5NdHk9nwcOENR0vm/fTeA26++YC+ixyLQIf
mOxr3ycsw504snc784uBiJPQstR59cmwYN9L/pDHY1GWDGtWSh8pMBw/IrU3gFgm
6or8vrqsBbcxLAf16dps8pZ3qxDaXrdH9Jo0yBpGjOTJSW51NxZiJS4y8MkAdKnj
6ScP2UWtdXds0MpfwFcQMFm3rYH3hcM6nTXjaSrt25N84dFK/e00uxycFo9PZX7L
ebZDBKB8dWembX/38PwwcvgUN8KeUSWobeZFwJTvUznCRDa+PTWMDhR768eC2RfS
HZkQ2dnA7wQd/We/OHDt7mKK+yBnJIqYONBdyGnPqKV45VubgWx87zQcGOL6FS0A
ubukuUhAFw5014kARtvdeihI/fltCmw9UTVwQQXwfdfRxlB+myT0p8KiUrA0fBbq
RxOhzSxmwTR8x6iSWaSTSCjCG/BQrniA41zsKk3uXLRr8pIJyGyVlu+Whmo5pRuG
IsHsDkF2ClFasQEr7NCjMQRIOidT39H0WXIpxhcJXMCQElGfVNdtX7jtEDZunxCk
lasJojTEK2jNB+BdhEl9SqfkGCMtU7eP5grAXWHStvykCrPJrbE2VvaeAo68h5EK
ysZTBMdTrJHeEfPhUW9rmeg6UtQkOWqnk9kP8Ig7MUNun0VgObfM6S+Vu6pJu28v
8ThWSrji5aCIOXun7T9byyOAmLvjIi0swKBMKKcu8J5dyt4jDDLACl177IrUppxR
1cWdMhyx8vKufMBhtBucyk4E6Pxz2SwNuikkm9oKA1WIgdwYGf1AqhoG0X8bBT92
sIw37D+HQDWGqAzTueqY/hQuuV/DrT8rrLF63kimWcYv32lFA6nfjw9f7ehF/pjG
+ZeE91VduencLDcuXOmiBCOBgUf0MESU7mSkGl8UXr52a7PddRq8/zmyswMT9+Hw
o65Z2X7EpQsaHveGnHVqT2zLkfoQjN7LF1YETz9rEGv98/3U/i2OaUmb7yNLfpxZ
FWuRuOo/KDrGT94vDd0My27P4hpAvKvOhS21Qm1ynyOhjUR+iu510Orr+F6ObibD
OTYsf1ICX4DDhfAVOHrergIkODkwLsHA9BvDliPmq03lA+2Wj0hK23LvMtm4prF2
4UVY2SLugdPum3QxHiXPfT3jd7Th1QrAyinhEmwiZ6XLcp6rsz6lWm7qa0v16HjQ
9xTXZtGgJnPG2EeBNNFWhmUxldgiM84515NQP+cRuv34EpXvVg01yO3jh6h8fgr/
ihCgTFeHnW38pMGSaKwKsdUe44PDTi8gOnOIB/NnmG4hvtQLgn9Ni/6IajS1QIdl
+hYOvM0o9kyjgyNs7CM6T79yDDVgmpjxjj5+fglt/YLfV2/+9BRw4gj6pcKAuk6E
w9G/HLRF8zhmA9//SUvTzX/zaHmClOcJpyKnio2FWgTVi3v+fDROd1SeAhMvAI4E
ZhoKyaLVT3ML2vPEVxl46gApiOmz3oZmt4eYpft31oWC5zdz0XSp/D8Hv6MCOXUM
`protect END_PROTECTED
