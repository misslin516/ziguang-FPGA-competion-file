`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k5aY3ZfrzirO4N89lZJ8vDRxeMGNCf7uM3GDd6h+iEu2N7c3HGcFy+st1GgHWyLa
WUHcqamIugcEbwXp1I4QaKXA3rnRcdsafz9vStlaNvdLtCEC0lU9ATDKC5XUjVmg
X3GaqqA7j0M4K08ZEixBvjy37EJEoDruCC0H2ZHJGhXDJZ7dOLNJU83EqzcsoA+W
SKhf4/c8Syq8CV0ilVmIgFxO/KZRYuUKS8K2yLYZqxw3OGYueJgrnpD9sVnCZC9o
xCeILaDKQnmQ6V5fjN9LiwXJDPDXV1Xidr5d0q1sYEytgux6wLEzMRCYeOZ4+Lhc
pJddcoQVfd8pUkHoh6LOy6GjQMSjcKtCHAO57iOPgk7U8ZWRbuHXxkGpw6JN+Nsl
DSgCf6rfOxCqM+INcAUpBFcE+mk+Gch1fsACv2Ztgyq2wpr6nnWG3mTuYe+9rseE
09XAAuCUm0OYTpNH7EFqH/5JaUnQIrwh+IuaJGIAwlKBjyC7lZUTXLfJ7EhyxkjC
68ko0ctzgJL0+wxv2Xn6EgrNL7QXv6wdxxOWQRwAcaPSe2Juk+Gr8dcMrL6DAUId
KyQfQAnOBS6yQ56TfeT19+NrLnoUgHc9CI7AUNBiSuViKK1T2r7Up/s7qJzUZhz2
bnlfQlshXkZGIn6X4BOM611LlDdEuReJaxHltAJRH8d5E6Mk+AKv9X/COZFCXNzC
8PVuSW6SLFR5g9coM0r2c8sLNLGqXvA6ZdtwTSACrddZjjgDJ7AZ1gpPyKQlg3pQ
/me9kErV5UVMkPu1MfxLNeNC7aXQxIBxVS2rDrSzeihRsypjo8nsIBjKBMRKW6zv
zvA8VoEhfe1N49epIOvelxJooXG/Xu6Uz0NJaIq4sY+bh6nY++xAHz2UYAtiKgVJ
FJemdjoup0MhP0/BQmFfV65BgacSO04FzdE18bejdghdvkdPEsHaQA/5KaJrpvEr
qhXX55BAO6uyXDATRvHs6TdMQhR/X6L3tcU9pQBFnOrIvpEThEwmgaYfePHOD7BS
qUUp6jfrGpX6BAT+DFn0RZ7YQNRUNe1RaoSEzpweGK+VYQU/s980NYcmD5FNR+0b
1mmofNFpcNGjLA0w2xNGu7VguhvNgHOCcrSaa62EMO0hoCP6hYSaVo1hk3QHENnn
YoStrcMbqDgorfadqsfCGU6AewUeUK4Uo+bI3sdYGEWeUyUGCoX80rvp6Jk+DzNy
+pZcuG0SpAgl33SqBwDgtKeKUlGaAi2axx2nZ/3BwYkfmpojLZC6NY6+Z9dSIiiS
CZXapLy4gX/kO4P/eTdw4uKPyIvGLTXXAU+ggRKuCcqD7iKF1jjNRH6ougaSbmYa
YQY51bLOAvwIefr5u5LUZcD8va8LtkUTYwsPAIsmOLNc2ZPD6UnJ33V1rfXfkPLq
iZ5vfKTXy7A817mOIg+lIGIhX4Zn0wRZN0UR3mtO3l7UA+IhcKcjVSuf7BErAf9L
KnazeYBojwX+3+IEHNX37o7ew4tSIdfUCk7JHFuR4abX6NLx5SbwXofL6aNzokJD
4JmAn0CfXuI9PfzcPHBhA5QoSehv09LbIGyPMDvOPdmyhzniA0ng1zVlaYtTB+JY
B/txAR8pNRTPXOgAusrDuUkXggjG6Kzz37azgqs5sbJeYH3W0dB9ZuWqW7l+lI7x
hi8D+eEIqJNKW4X2b3/qg9BE8s21QHCrwMWK2rv7axBizadngKvOIrn9JcAvrCVC
wKqwm4G94Gqz01rnzL2ahA==
`protect END_PROTECTED
