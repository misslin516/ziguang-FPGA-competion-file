`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TdVaIMddAVDq7+RL1ildZTXrgQw7KWSH2trnWyEi1NtSO07hnqFCiMFSRIKYUp4P
QE4UVsbX9s8rTDKvoklu6JPvPkiFoJtoMW297Ota0Nc57XTvvhOvypg+OlEJJO+Y
YuKEUo2VuaQhmXrNlrssHbkFaCa+4KVEnO3GkzJ0fCT1LMMqbx8L+CgPb7AMHIgP
HK5llVbqF1pQ0GxMe7El5lD40NKp788fIl0GsbIdyrxRichnh3kznDnPyrBY3uFv
yvYU3JWDBYSHVYsAClAu+9an24sjmVLJUjyh5qeFI/P5/XlVmM0H4IPkxpN8nHWr
HyrcfFGPSomduBZFP5zIHhA0CPBQ0TWW+0Wm6pabzs2kKNpsEiZbS0B+Ej7/gMwt
ziGBMiaS6tWp8FTYw9Dap8QTms37mYEAnUCCz1Rfo73GFGmyZZTe5A0y+1GaU2C2
R0mnVzE89lfI+kWnFH3f+Z2OCiH5iGV6xYWgnz+D/anj9gecMf13wPUGzfSc/HKB
YTuVmwOuIvGvHqUiyC1061OQdhnUr44c2sOhGnECIXuJbPPtPgXEh+z3bQbrEfL2
8/lhS/xYkZF06i5MmW+OSBmIJzGXdo7poNxpL+T//7DGWOXx2mpZAfg9KCsTya+y
DxIlgDf5Cx7iAI/MHxy0o53mZtzyIDlZEWONDVt6xr+pNCfbqS5oQH8EKV/A3yEd
GFw5NeBjawtB3GPpth8VjfA3zZ/zLbu0ceL7lu/3XH4=
`protect END_PROTECTED
