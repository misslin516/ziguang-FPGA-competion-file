`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCSRgHytDVLv+nf096O+LHpkPsUgWwhPBqIV0R3xQDsd2g5NjH4BwtbjjObMPexg
Ig5Zi3vrM00wbcczkNmXd83X1aR1319oJWShoE9ulSJZWhdZxnHldlr48Zxrs+eI
loOBON2N7aVIIuLPbky9JQbXtFKuAfw54/NkLz33SeDkJH/Cy6wDMIFdRuN5mjBW
t+TBn+O3Ip0SXUMULakeg7SbJ7IYnvhDJOiQYMirSGT+ZE3hQm1chHiCi43GR4+a
GPhQmcJHzb/Bkm4MzPe07WORVpBkeEwQIBCetuJj9MfkRbJwc79LMmMSEFexyxZP
FipeMIyP0qSYFfncDPBFf58uL4gb1IhjQcJH3jIAIXO9Lf7nJqEP8Y0YVMgH+zlw
+wrwFOQ3E0jK4OBfjtZTHKwK8sSiVfhBe+STEA0elHS1urgYfL991B8ExIfRHIjn
q9cFiM7tnEBs9m8LFXTw5nVUdakDAG1QsNt6fmFckcpGoIEu0OyZF1mhesOf1mZK
iqDVuUZbN29QW3jbWgau1zHp+mNHOHzRJYtXupIwPI/9il3Osd7Gph2LWxKOr3n7
O73MObbTX2aI/vS6r2JF1/+jB7Tvw7bUJ69ON1DbQMerEd5kSURAdnVX1RebaGFS
59KKFUl3VQaFivYTxiweYcOjXeqX+5VKY2w38qkd9qilYKs+cv0hRlUHcOWRTxtr
yyjkRMoeTnLwBy7+wN4613jCuEQAqs7qf+6z7SriHH342C8zMkwUTe8/8WaigJux
pQYdjQbm9SWQ/cNI0yVVrKqhycXS9o5GULblZKhBpEW/0b/s14X7gYX+3wuac59I
UEQGXIsLNzlwQT3Oqsdc2ujI15OBqZjWmr2tAVXgsgAs9PUk+Zd/YHCRQcOP4I4E
ZzclUhO5c8upvLoFkAucWAXh89fJ+tPXWXQMSdfnCv983g1h61nxq1ShOMNTYfSl
km1oV0rHqwDP5RUoM1p+XqAPkbdgbPbjaQ7sQxG7AtaV1ksBnzaJEGV1vQ3R7iQF
IRbX5DcHCxz8sp6B0j9gSPEEuaI6WB55soTtzlIwfAQFvHZUI/tASGpK1IlfyuR+
Js0p0vw3qy2IvUgtb/bkiLYjcoRwwcO7TU1KDxsufsHhly7pc/nQh4hHQN1Ud0cm
nPtikuhPQyKHJn3oCmQckNzdUIBm494gUDN7WCcnJqNEPXs/MPTFcyFjsawug9mf
CPWU6k5HkIEmNWRMbJ02Pwiz+qrd0o/Z1yusLyAfd8YJECcuXykTne6BxEit5xlq
TPWjWpceCBHLOKCVOHEOu9SeH4Kh/LAF3qDgXxVZNKA=
`protect END_PROTECTED
