`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6HbjkteVLJdgO4Wm3A3aEPZAQWQRTUsgYCMLsdovuyiOJTC+ERLEw6hoAQZGTwq
NJ4b6Wy3PAux1YOFR8jpwGEKce0x/6og7/1ol6hag2SqmxIoz4HnUCy39yDbhYxJ
ihjHex/bGdZccacRBXXinPK3eT25PiHni0ano2ePihvw3o5LuHN2GnmGH3ipMZ1B
yCgdSmgaW6/MUg2lo91H7QDJujkevfdDJdasJux5scktIkstIgktswueBxKZZYol
n5cNSoMA/Sj9ZJVPnD8pSxJ7f9yyX9mrDG2Kor2BjWexdjY8vr6tU4xan4vscKLL
dLfQkdadAj8ZKQKCGhTjiRdzoFQQFBIf5EukDaCUIuhBW/v9mGALDKg18lbZkSSI
veZiUnKy7r/SJZluD8H06BPpxzS7PdUL/bFkX2yqYGlIqSYIGKdEG2Z6Sx9e2612
ZzDLjPKgISHOQoXEmGP7c6oev7amMbM6hZzXNta47t1pWtU4b2gx0rLFWq+ddQ7j
WAulfW2hT3NJFS0F1d2TUNACWrffL94+MXBbC0Xe0UWGOyJEGdfs4NUdcTreuCHO
c8bv9MfSN0UZeRGhHzADOccgZ4Ch4tBRYWetksYvaIe3xlA+t4NpK7CxibtzUZU5
CJYciKZPSI21wz7S7BZikuUl0V1139WGZr0wL9F5zyxZ+pa6zP3oX3qCIjmzK8it
So5/o9F31CpUl4EECiauHVifdWV1LpL9A6wzw9eIBHMYwnsqlL8hL+Y+xqJsmKGX
vfDlC8tjClnIpc73ZSXFS2wo3HyfHW9vdSFnP8wKoqeUeKP4Cp2q7SpvZwJqYX6z
pUW7q12ELWkhxtCfypucI/OMsP/PaXupKtCY6IUCI1PYUUIV2S2AEZYT3BAGx0WN
AoMr43rLkYCexkMqb/58Wxbn/mGWGMZeA9v+V7AeCxOmMBmCO5QTvGyD8biRpooH
NtRJaL80hv/ZdPdJ4m8P2wMdiUl+0tHd/pw/ex/kIvE8t2Kkt8l7b/RuXBqnz63B
oZRINzQFlE6gtwvGSxx1He0aj35uz6G2F78yt09uZ0Zq/x4ZlY1bHQ8hWXGBSAbn
nVU2OnDuWKaoluTx5PAt63DiCwXIMXNhl9Fq7wxD0F80M62j5eD2YFn3JMw9gu98
aJjlNizLxD5CMnrvFFEU2n9C4UuduLiakgpPtXhrC+B8fnAW76rJC+XqLGPrNq/a
C80hq8yccEQzuykra4y4QV+NxRVS5KVWi5Pem/+D3WxR3294fscjbqlrtulOsDx3
AZ4LQpGnXjtUW97TvxrQ8unQtYgUeARIfqzxfGB6X/uT+935QAHCvptWqG/Zz/e1
3gio0vaA7uYplgFmRpIHIluPGwpNv5Btl9y+JRgEPHJY8t8CD3QizwNcN3uvjNh7
PKZgNYMJ0ng7sPPdTY7JkI6dZMMJAlFgzvIfcHvYAAY=
`protect END_PROTECTED
