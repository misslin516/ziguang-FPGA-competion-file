`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdv27DR+Iol0/+BqPnfzQkYZkKauVbFOPVDfWxY8wV6+MOPzSlJsddPCKmVW6fHW
RhrlJKDhBxwAPpW3C4sko4PirTfdhNTc1on3TPiVBDoeeipmaXL+5KHOuvsDN5Qo
6t/bGKqIAR6c0vPa1Emdi1Klvnj/hPXnnfZhGjW7KEHNFvfxxOB83vCfzErposX4
27zgfIyEHrm7D/QwoXeDXh0P7NSppjIY/OzFHbuQQj+RqpEovPIpq2vZUiK0A0YH
THekKEXQEXRXN4Z/00gqx3Gx3qV8pst0BFIepvjFo16DtVBSQehf5qSeYM+VYT+z
v/lLnc6xxmvSNmPGFJZZyDiL2eBKyznqEyVesbDFLVmnHv+r30rm13J69D52ujyr
eJBc3LvpVF21JcfCLbvLa8IceJzpsj/kBjxIi6j8mLvPLen50TMwmXKx5TdbTsAR
/SEVGvtkvFi7t3h8B75iDMRaku4QFABGgS62MPbc//Rs4Y+BetWB8EQkURJbk238
qpO+8f2lZjXfvdYD2qJfASzOt7amsHwShAQ+4/RWyjVMXsLYrL7k4kACZQR5MKZm
+VXsR1MFcHIGZ4qQ5rZYhQvNjzZ6HzSD9Odnxf8HSLz+riwdCdWxMUvcnPH01cFo
5p2F9JlRdFN4C8IFh/764FmaV9g3SnsShm5DJlxb9NgZVpO5ttyAUFEYjuIRXAes
TjgA1F26rmvPTN/t1TGk/QpRCi/S9hKc2HWBXt+RNFCG6E66GmoQAicaKl4h1D9H
27TmjeOU0TAwueUtBhxBxJqRVggP+W9zmkZjfOOF2IrUBzqLowffHBtpc66309dY
cSpl14Ht8a6LjVT8LH2biYA6OJpr9/AnHDMxI3dIHmRIRel+HI/rBV0y5YKAliSa
0IjbWoRe7/XhbzrOUsCmF9QG1s6IzqtE/YtlOPkWtr1W4IphJDOv78MortBIydrF
rgugzoyLDmJf133uSEVKjSPUnk0Ixy7OGHn89yfcjIRzOMf4ZYfdEobW3UX4Nlsk
KB8MqnZn6ISCjm566EEsL0FdCLVrgCKBKzGOrmBHkAQsH2u5L0y9mw5biNxdxbpd
m7Gxuhrzzw7XiO8C2BUePm/LWdZt+3hy+jZq3ngadNCVIGLKTkH6fzokOUVry+5y
WupKySCSuBbYkAXIEChMjv7ih4IlRa/9CnNA7EeNryTikTYBeqZ1U6ZPnyzTOwhU
yWcqAC6Im7rIa5P59kE3BhLwVlK9xO0ZSoXNNbqkXU92woaBSBd69CokKql19nuo
MjryyfXYWD6+DdINgS128MkhflOl2p731tYAdRvARwXCVUKU00l2KhCL/rmi9mth
ehN7rKKAE7zJ0OqC5vt+B2LjAu5MgHO2QSmU3fusfQ+WL2oxLFGo57OWdy7XSyef
KMHNxs66CGT7KIfMWJOt70J1mH1gBgxNpD1c8AVDTaqo7sH1s9dEpa3M0j30/r5+
/dLqbIwZ418LEX+9ek95c0Zw3hOYSkQoqUx+uI9/ZDlg58HfE1jDhqt8UdXcN9ki
xIJVzvnVRm8KXBcYB/qC0yK/DIWa/WGOogHqI55nOScueIPCISSZJAXznJ6cTQh2
1r0rfKB5wne30C80UIgABBc+OxeJa2AvRYR72pmdyZc+X7kPdeYpdVec04U6gNP/
LirONs5U42fC25B/1gZFsXXrrvrStOiYMKjppqzoWmnrx2xBjGw0FXfe02uWqkxH
bLp26Uk0Hj4b0e8HqbUzyE6/7CCap4YBUSMd/neN7ogKlmDBljAjMPMYRn92oX+a
xPjxabLhOh23EFuIZzmZCUFssL1V3Mos45KOLOWS/VkMQxO8JvgweXCdU7b9SGbe
7qBiaAx/K59lVh3/AxutD+TbMQShjH4d/JqlVOCwyG4grbTySgp/D9LlowolwZ/x
b+j+ObXMJkD6O/W7orUqopB7UCLN6fEYgQ+Lkutc8DQzMlDcvgdXXbrzjvwSoePu
E95t6pU2tDXz4YZrqjswGxfo4Eatx5p2cBpj+T9ES1pt2mG/mWyOoCDi3bFxCMfY
HPDQ5/9BcEW+EruDsrPMZqgU7bE7ZF3OObKLeAjcvA3ZtDKZq2/FvrwdhHKHgwO2
GtEr9V4/CroCqbsbr5Hw+EJi9y3D755bayDrMFVDi3xIMxh0JwUQzzjNGFhXzXFe
f91INLUHdqY22XuabiS1t7MX4dwl/JVB4lcwrMZhYC6vLSGMQO4jIpHXMohwIQ3e
n7/lHZwsMs49lC0erxp4zvqvNVwCn6fMpGEZZwE9Glq2SicDgeRJPU6B8TtlRLLo
l/q9j9TKOm+MRDiVUAAZOud27RA+oRW9pNuVrog2VzXP33JrDH04w0O+T63BNoC4
aAi4bIo7TcLhjHfCmeSqKZG77KUdrb6S7t6wOaApLDcP/CxRWu8BFIC4wMETLZyN
xEBWRuaWFHyJcvZzPmdvxv/qEARTnP+QKy1Larwv4U+CvcDAr+3fnFtclU61FqCk
ghXJQQMGMPYNn5sq/vERL3+eWgeIO54D2jv1sVhmgn9LrGVxU8p8qITvzWpEeiqQ
l7ggnJZTpzTrH8bMIZhnyr68NzRaDD86vGWzKnfyeEo3mSCuf5NVfe5V+gGwUxSa
OSnFV2ZnWvzGAM7/t2ZaM7aZFKvkuz6j20WpKW1mfkXibc4rDE8u5fQYiacqAFD1
i1mbX92VFjAC9kaLQ9rShNG9HHMl5fQgXW8xE+7T24rF5p9AoZWb5hI+xrd5xtpk
wFoiS54PUt1yCDPRS7wounJfmbNW0sGJ1h6p2isBB3lkE66aGPeDKO+I1KG2IZZZ
YVnxmXhd59JBIYvZMOpnxOQ85iv0vZ+R16jxWsbzCdYHwJsnLxztPFSy/kBP9VBP
uv3IXqEBxvGT8QjNI2+zo1W7g1U4o9HC9n2yh2ymykUOnsfS3aQZy/4Oz05XtBi7
zTOc/ryWjSx4bmuQXVWdeLxnTa5LflsyRn9J8IHF6glN7rIjgPb0RaHrMoqGxBAV
bdTRwv0X91sRR7ZTu6xV5ecjrCoHTEf88iDjurCAENWBJkBD2U+G4Ps9E1TqSre3
UFAqi1bM+QCYdJLhOvrAl4KLTZ9Qh/HgQ6uj8ai7zAsjCmp2z9gY4ouuqFzc+zjK
eEtll8CCKyvVr3qjovrLq/IFlbzRECPFRZu3EgqfpnivjIJA2LfhEea8ibb4UQBC
ei6Y/J1ziQtR86m/RQJgakFU8S9X6NBaO5ke7kuWRLnfiUx2ApDWCotDUGC6H9BU
KpppzWBlDQW4bfjDG06XijvZMVKYZ7eDaEYKypb1tEGuN291w3UGfqyQj0mdeJ87
DQI+SakqB4rx5IfGGuEIe7bl2Fvn87Ehz7ZUQWEVQUGHl6fdWzoU05ZTKgNADn+P
Vo9RaTzEkuLRKE19cfm1kBQK8XV6jFTBQjFE0ILKXrhdkORM4eXcTgh75Mc6COkr
MCWku5lnhTl4tx6HpAZWsXS9tDKvnABU5gFnaGmCcz3N9+LxXAzq+1LTsWZboMB8
mJo1Kec8AOqlxG8QWLfdoGhHo5ocrv08l8aWszUA6QvgTMpb/MXmB8hU0ivzhUe4
47Zch/+l8M0yMexCK7tijW9Cbmo6dmwktZj3cuabuiZqAAcxlCEUMiY5oVEV79u/
O5EN27ldewqd9Fcrc1zm5Ac7dw2J/ObKSSkJyXhQB/0uRi97AXkSc/tyXRvrJoG3
t9uKmuoNzJLzZIgaZw+Xnjpa4/buwDY8wz0gdhnbZKrsZZoB/W6ZBcbtEMveWTUZ
Lq7O6g71CVgJx7w2Ok/XRG8Mb8ckeiVX01yOcJpF+0rmWdZq/7dt+GD6k5GI+hIP
7+1xAZGCR8+qmFrC6dbqxte6EfMMMewkUy11+8iRy/hl/Mag5A4Y9525jZS98r6J
y0srHsaiOKZbSPqkP2urQuPh0wsu46tZJ7zPwdKJwe0CTlHXzQcMP8wk1sz4VxQ2
XxP1XR8rwzB7DYTMuttGDe5o9tfmi1IpEsHq7NopYr46GDtqDw3sM0Al6NoQQW8w
avmUHj49Hd/8VEQW7V+eBTs6p3bBovvbBT5yq7tet3JN5Vx790pGvoLz1LgBL+nb
W8/O+Ad8heNY/5huSjBlJ5y1jip/yNHxQvrytFzl72D9tijOEMd6Y8AXKOiCSnDz
`protect END_PROTECTED
