`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ygCUlYfGC3jtkG/86RTThL5NiIB664Z2bifAEsc8hDHUzAX1ZNhgy1wgjPg8vkLb
3RCMnY/ZXY3rzH+5lmVXNt++ghzhpbq8LNRBv5A2r6jcppSy/1x0W77kejUkVLXc
DIIE+/F4+FT+3tdM368G+OWNuIUZazSHYApxyfAtSh+Yiji0D8neBEw4wE3lzYDw
eUeRpOTFlYjDFrzmDWqXWZzdbDkF4lNBfCAl7ZxwoVRIDhMEK1ObfgWcWqfRsRRT
7auUasc2r/jfIQU/4xfjDQOsBHewrXnut4sf3uXiDm7oDpXQFo59m9lDsgxAhIiI
TKjiFKaJJe2m31erI3Ab/6x4gDRhJ10uh+zjEtyC5cNaf6vHDNkbDvYqlSMcewhA
1+DiSSXGZK9iBtnZO5qEV2pZglIo7FmzJu4Tfa1nQsW1RK66SSMfS6LlcGBUqqSs
hrdXqEfiH+PaKPt07aiaACmjQYKYXoVvp8gHsrJu74aTk4YnXZ5RTgteH9obOYjA
OqOOI7khEur+cv69HaRurkc/PGx1Wolb7O8GhTT3zSMaLpzy5KbMiN4b2fyASQMK
kfZeqgM0GWQN8EPRh4ktQ4yN4/GJ5AkWUzKlIEleIJAI3l+//2smPxB3jRRf8hi+
ZsTTp1A8aPz2QGxFAF1kG30mUixofC5Ofjpz1BHEzTgp5YjASOaPofC8L7dhkHS8
9RDQsD2mPPEpyxbp3+cXOB26rfErdgiBlaRNim04f4K04x9MH9+IFG9bxjAPlV2j
qb3QkKN2rYC+avCyZQ475kpcSIwC9OkXEFE9O0Wt/mL2a8ayNMubmh+4hpULfFTp
EH0qiRzERDb9jlQT5NRJMX0P32vKpWwGRRej0TXer8NFeV2g27/YegzJn1vWm5At
BlyNChifxZ99ebdlT/kBX46oZiHEpAytlLTz4Qh+9VxftoJSDXirCWku0Kr5BBXM
2Bh10laJbrIyxPt7qobHTfy6FJoNB8ZHi4A3gCVlHwmlaHy5mudxOhu5FPUldFAK
RRPXHFz9n1cDWAkvQANv11MEX2gz6G1thhMxMRwRg0Zaac4wyOYWK0s+3+fl1ZVq
LvDaWZyyB6MtIYbengZNgHFzSFV6+DrdiOhSG0vRj1miqWXGewg2Wd8YgbluIJWh
cTWDW1WCJpjS2ua/Gz5xbD8aeBpW/z7ufdmuoMRa89kE+g40K26q2xHf1gcg4EmQ
35YJZ83N4iAA4PvkdywkLlaezJIErRIqO7I+oSl537j+gBdVg8csQHmbfdaTl2En
VQ302t4Mooj6ZeyoMPGl1DsO2B10f9jelNj40R2Ftlb5o1zSBYA08NZ0vefNXhZo
J5llZrmaPctSukzsHeaIKyzngb42s2XeR2vo2ATajWwu5xA3ImXxiAm/1ZC0dzWm
E3qUrjOMNoU9fdBxLkXBYJ77ofP2U6YlKaAPzn5TePTmcV/Jp5ipx3c+R6AI+ZCL
EJP2pZTRI54RORYj6lDYHIFSQnaIxI5ZZdOrHrfDf1stOnfwqqbKb1ZH/7K9PM0X
YnAMZDRu44uYX3SnlK6JF6o/y1EKhLb+hv6ij084Ej9NBrPFhkMeYH4GdHuOaOI3
KWVlUat4+MLoVp5bcRVsmo/Jc7rzE4ni7DvIJQZqxL/chi1nVPXIMHPk2DQSPHZg
KVRm2kNxypt2urDEkXSyaKJx1RU4v6j29BNmw4hImbCZTZ/6S04+ZGI5tN1+eLJo
K4sMv6Q84eqiRYwuEuFP6KsFVq/fTERlaTePz7gACjFUOpKw2fg1O2L1JhVou69+
SJOOqgsqK7BhXX607K4FyRUrMljmYxlRGmBTK4Z/B8SjUXvNLBWo6hstDrAYzfvr
wwGH/a0OeROZ0GeCcxntEchkcDDTEu6ZEKEb7NYEXPgoGpfasnagWizzO3REnTcW
tUopjn+aSxPGHU3T1b5KZa+Xoxys5Rx2oU9Troyt/nOLLE8yod32lsuwSX3mkiHs
amL2VG/Uvezh7njMQKDjrbtLNropoxGQyBSOVULlJnOYB5XpJqlaqf+xtY+tpaPv
kSFbNvqRmB5Mzek+3aqACBrBbnVE96yWzks7Z/c/zRLMn/m97Hgy+tCLgb1jEM77
5m60zRW0+KXTndKBybnTaMjosL0WD8SmFxSuFnaax7ZnRuQsgYHTbliPUgkiQFt6
20+rOtGALI7hRmewk7fWcgpGN4FHzybtepg2n0mDXq/H9w2+hahJoGk+GY5kLZer
wo2qXNYH4tbbRupqnEWBM+/0zOnbMenlTq2cnyfaefLT9F0k3uNN+eAQxUkhj8k+
qZuoWFo9Fl4A1LKFgNQ4voUOmAPVQ4UZ7cmUUmkRSU8XvrKP/sYjgM7Ln9WwT/li
As7+Tq9dNL7sO1/OlwmXhFLBSkgCJwgOCOOkBCURixe/zyrpNXnlw/p5EkMd/ho/
dEEGwj3pXXO/gtr2OpZihJBADAE/kfgVx6eBvpbKb8v2HNBg973YZHnOurrwuI7R
4qJo5GXiZLs8RcDP2znUpj2gG8FJuo3Uc2b4DRJuWosmWSfTUYHG83YmrSW6itpk
P3BX+ITA+YwGPdmfLCaCwUCBmA02MCou6k1ziSsN9Sqj1BUz+otQjbkZyTfvrUcJ
`protect END_PROTECTED
