`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pp114alVrPd3YktSVpbupJFU2OWvAR70eb7bj4kBByWPfeGLc0ohnJvAbbHKoQEY
cAApU+Q8Bvs5bIHR0yplemDxpre3BYCWXwK4dKcSvZ2+c9KrOE/gcDbOwf4FRcnY
EEL8QU+crBMGPwldoFOtQ63eNFjbILPESWsg3CWF3Flzq101b49qnsVxpfLKo8on
DEw5K3iBxW3nkHiDTAhanjjWcqxvx40Rm+FSF21teHUzh8fNywHtpOqY714hvqyA
2vc1vhtJyYtsfOaGf3ZGOJiQliY6VlgV39uwoEskrAoLRrIeLWuvDaEUINNI4Oj8
IKYTtg06rIXqho58bu0qUO8pEgmJD2VW+X5pPitCez2HPJMlaizrv9+cH4A5MGxg
lVY4IYggzdAL1OMrMpHutho0vEf70aSDSCcv08jOThMQz44Q4u7eKcLcQ9KmoQlg
61YpdfW09NQ69YwheSSBrdEy++tz2wls2aE6ztV9A0vxrIEAZUKPPddBsYFU8noB
7yrELETONoPsxGCLVmwJc9Ul0oWCeupPrOmhStUM/HTwCZ9cwwF6ohv2gI3m8ueO
odz0b+bA7NOqC7zMhC9hXLqVnjc8QqnOaPueR4W+5Bw/MImPxvmWX/UDDWgXfjat
niLeB9EJ0CjMeUzeVmWm8S7+0xsRWGc67qprax3kSjVCHxiWTY3ajlUMsAs8ULH2
qY6WgoM9LzIO2l9ZBEKpAlDAhLTlcOsxdf4Avbv8Og7jD2deDwoJMpElpwYObrRa
s7Ngo6RosaFJNZ9LB9easqhGc2VJay52sZWkfpXLnXTPHXGp3N7kpzvYv5PWbeUV
KL5H0W0dhja0LrLegWmVbGWE4v7hfcswfBRS6CzlW2ETbxbzakI43WMSaxXMrKE5
9dsdaXIvh3CT8GjWobUguOsP/zvdByflCZCvJ9P0clxQpSCcAvnfa/mjBnuFBY4L
gj0SeUHe1xsjn9yfF1Uvn9vqiCBNhtRp1Xk1o9a3egzFoSS3DF2SNZPQA35gNqDO
aWezu/3WFKQW1fngrBjwwFICIVl6c3XrSBnCoTk/byu5WnLFAzSucu8+CLRneULe
OQMYMeWtbUiQdAXAym79nthCt8B1Lcuv03+ee1Wz81CcSI+azjnvs0bE/DeWaUjo
LGydBM1L6ac3lzYL9480IS3dTSti6Fb0YrCPvvmB/AhV4pU0AhcUWsOANUbTkc6C
WMn/l//23OoHNDP+89unncsmLNyOyy6oe1TM7AoaQV6sLo85GC4w479NEP1/7vti
KhCDVY/AX5XSXsoTKeeBw/E1JOLpO64weXl8133HKHHIh0nKYJBZc/lZDIeb+r6a
f4ag5FyxcRUQZjug5SV9jXwkiE7Lq+wg220iZu8o5mLCPmLahxwSmB1QOHd0Ucqj
Z6FALl6exjI8g8nLLguRFlMFHWi8Hn+g8qslob2W0MIF6a/Vqjfuzc22OxZm/89I
9MrE9ECyiAZkzD2SEbMabA9UT8uFwMx6AyrAQ/noDmYw5c338xcqh4djN5u1Yd3w
pViDsXuy3CKTLVcAaGXiqdon+4KklqYJVoSb70aQ5fj6Xvd85ddWiHeCot/kRz2P
5B8MKJRX+ValDjS7eHyjWdGlghnDM4VSds/6ocPcU5Z8QNiY6Y8OxKHCKhI1dfJ9
uDrRcvge9Vz5VfOQOwYe2aHkmHC+rweZu5J+D1XGRfHf3GFEmlnbks2ZbmbUS9Qz
YiPGOpu/pdTHO0FxGGFJz3APmIv2OT/dDYRt58C7bWkqn1+mUqZfKvxaRmIWVBpE
q3GuVitld7oJwXpEen+b9AB23Sd7b0W5EVOhI6rwubkfd8hQFVsrerf9SFN6Zu4S
5LYYySWhcnrnIBRTupydwtYNyhbScFSCtrgcciqC4CewHOFBFiGHrrJAxb63eNWX
GgjqRE58guxbdNidpU7xAbE4sXSubzggJclbmtBfmrFDAy3VM6y9e5bB3nDKW0ZU
fxQzCBsPqn2nr0iKy7GL7fAhUjVRxKN8PSbQK13a7EnIV8wN48JeTTuZFRnNdj/r
iSg1xJcHv/9OrvLJ9/v2LlxNMX0vMIEg1Hgmme8MzcLUfYB5SnnIC33N7Q+nEc/B
YVAtU2zGlTFUzImmLRxyhQmH+SE3BBnwfPkmgRYAqB7K3Qk69gqXvwB/vse6d4jw
HMkPxVfHhhorOBdmJKXGC7srzdQWLCYMlFUF1ae5OzcfTLmWJ7mwU/XzSoe0/w5I
qhXSkJnkZ86eG+5jZ5X/+AKthh2W+eelmEfpv1mN03tMRvs9gcsq6kqBUUeG/uUY
zGSHIOxQR/STtvrXpH+fxkLQQlXIaxQOUKKXI3dd8cEjOl5sFNCPEBMG9N93GSxf
1Qspu5+IkfLKD2D+BIzBAR51QJ1QstWy5W7iy3KV/e+I4uurY9CGQfjl7V0VeZxn
lZ7ZucN/KY1D+vfyyOwiPIva8aJISTNv3TCS3MAgwzlmNtamYyS1JQpQQXhOKd56
HrLFOEmn0yV28AmIzJO6vE8ZrPNi/9yL0/NuphpNIcFMnOMKT7lO4YNwgQA/J0Zm
fO8TSk07rBS9fxq0CJuW8l3AOIfL9YX+4nm0hogA0EfJbxQcEhO1x0tnAcwsLhj/
3c3OY4TOvyzDAqnalvP5r7WjGBYo4kOTxDdMCk1heCU88zNwbuUWwccWmJy6Cu5K
en8DD8WFMp2GhGo5SaWQf2ZQxDCqfN/0zfM9EQ0k+WzvF+xrpZOhKA5+15YS4l5+
ZY5DGTnLisQXbRRAmUxULfB6Kl8S9rLRwBoVHvP4Zg61ECHzeWDKxJK49M9iisR+
i9mZyknGT9s2ooFVXwrFzcr/WaqqpqUVjktVHKatunCn7sduwmQBc4p+Q1ghJOVi
`protect END_PROTECTED
