`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOKJf0Q+aujp4ig8cr88wf5BdoxoNxonDr2yyrrtBDwjSh4T1krIGhCooZpUB5xD
dwG8FpR2X5GfQXwkJn3SbxBKNoO7DsCS8PpeUw15lxJJSZHaI+9GGrHkF6GksEed
s/X3QGI9uh4+oXOS6CT9JEfCq90ZKhZJZwXS3l4g+cnftSXjUkDsD+/UDtDOVEvf
t2Zp0NxwJ0FGeC17yVQaxCJ8dmsqeGdDLfqZ7ePkWlv32+AFknvZqCB4wMy5V8w6
dgS8zBJWok5Hh9xV6Li3OvxjqUtLWwmbzyPwWRlPYjN2kqfHtEV7V//x0aq5QbzG
R8OjCFhuunuDlGyTKXsKBjzxFuMn5taIbNSjYyN7gB8GIdpgNv5RXCGuz2wHvyDf
DE66IWa0PXphSyQd71rq94iZImQIh2GRkJCrp50ltPxTeA9tvOPGEo0kriGjqzzQ
2uiR6JJwTGzku4JQKHEXq+fe1FX5bge/mg7LxpZQzzBhfGAXjjK1pXgdZnwtC8IZ
DPmxHQoxj1zR/R2LIq0nxWtJ+GO/HxGEkI9u21wC9wiooB1T5KaRS9e9sa6cFF/T
uUHlW3yPLfj3qZf+lywzS8rUHnDWLkLLJbhaOYCczk0e6LmOYwPwD7ovwHShWr2S
5NyZ/XmyU0015O4YAn5YXNLEK/YTt9+ATpfklBOD5pG9Gbolru0uTacK9X6v7Ybz
HV+YLKtnJxnZJP+Q9OaWmEkaRG/Ssc2IqWn91aGC4NEsdfH7SjR+qJRF/yljBkYw
ieLyfvqh8hvn+akWl6IWG5eMyUBkw06JOu2O2881sDpjSdJeyN1bzgDWgjU4iShT
oueRVhs6LNKLSwQM0If0otyCZVrlmQcokdAbyDXDGfHnzx5mz6zvGi3VK3PxXgVv
W0jTUXdfBB2QCoNGY0LYRdu3nlZ2WQaN6yQGcRt/K6o5Qy8KRVZtgir+wIJZZovr
gRA7euSr6S6c8ypvYtyNgI8X+7BBqi00/Z+3IE8umfqzd0zdKvNffMKJnpvBq+vV
ezykC0U7EBq5EDqd8fSNz8ukUm8qo/IMyPhO4qwUUnt8VdKtJlMl3dd5DkRjbXp6
3RghFrfZnXSiTkJj2AzHZVMEChSDgSZGiCWc5bAv7cI8Ln67LFfeTT5JbmYej3D7
DQjtjymeZiiIFWQj1XyiVzNiSujDObS8qpt1i8/cXCtjH7UbEBaBdGZGP+13yLQH
fph/Gn82oMgyOpjseou2i4a8z1yr8NT+TaEcr6/jNWAuEwuuuLxRN8u6po0GZUAK
tBRSe3VSx97a6Rhif2GUoxzwIl4OVt6H4xGtBTfq1eSmFiXx0wtI1y8601dBjhwo
8osTvIvCn7MO2tec2Q3Zcy3k+5K/QdWrTSaBgtCCJWQzqa1Sr1j+uJjRiSdVA39d
x1abAMv/IrOgE1hYtRNsYUFOIyVNWacQnSlzc5N0KGW4NLQtLW5Cf+qrw3wwy9xj
GwYs+bIGXqIJot5l9cLdOBMxloP7A9QZTOUlwWOgs1XRshWTU/zdO6vhQzHOEj+f
WGlMw4SkgJDR7+mC6JiZ/AgLPoRJ/BFYPt4N7PhrmfQhhDTIINcVO74/onf9rnbW
Xyof0Q7lql2Xmhkz4mp7KoyeNZoZPlImKV1t7I/7+Z1J87iiLDXKRgLtGxtPMpuI
M25ClQk6Pzoh3kTutW6kecBlyE+N15Sf674rGYG8RY0YQuVhxuF6+TuTr+RRPUyW
J8PXelcTQYkYF2C9COf9vfzNp2prMGJq/6SYBVelc5Bz9+fgz7E+KW9qM9T2S7GV
SYdqlahoM2JxbaoqGmlH/H3hlnJcrdpg/h7xLu7BEfX7pegrvoGlRVqKWZ9GIICd
hpW0vvQFSuEJufTHn3IUqKPaindYBMh6hs8bEaJASmze1dX90Ebp/UmIq4C/N9eO
ShC2NV0ck4iXZo9oRQgqcnslxTO1T7qMrR3A+VakvGHnmKMH+N3Q5fEb5+w9ohBB
8J32vnvWxjNXM3HfDu1dT3sEEAMzazfU8WYiQKbPEH6kMJfOiM9Urr05jU0JBotk
X+dNJEAcIlmhFC/0HUXjEI3xrr9iZ9g94UzZT3kPQzdIhEsbeKkVxIN9+QroPTIS
WZxRVY5utwa4GsTYHHadOG0w/qDKIHntCjb6W9Sbh5YQFpRpKHDnJVL2Wy6nKNP7
yNHnZyZNTTI17f+EkX5QnXBA4OCVKf8ePjviUzp5XD7yDbAEZMX9erZsv6uuP7dq
8nih0egN8+zl9rV61ohtwUF1PQgf2Yv0ifvUFhFtp37eykYKrW46nXNI89EpiJ4U
3qOf50i46j+vzBjcalRfGu/xGvrdxUnkBllM+kNmOqs09QVPKdxhQiGd4BAyUQqt
owalp3t6ESaf4IXE6Qi4VK5xAimjnifDLW7NZo51/gH6wSe7wsWZ/YAQeSH4Civv
yG4Mb4I9UEi5zBXmhmKblFbcDgJfhokp2Xl3yzzqmtMqP2//e6CF/qS0LUhsCBNd
bTHiJRShgMZyHDr6/G6cq4Wk10oOJN5yiLyRZa2Al9UUYggUwQX2nOx4vsxhXnr5
6C4PHxJIZRg8wH5l+trVZx68gP4gVF+eLqYO54c1wqhQjO3P6Yxr0nyBZmbE1zPR
U7KQ1tRs1ZkxvGQkqv6uEA==
`protect END_PROTECTED
