`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xxf0JTgb3YriEfgvsxC5rOIeUEh11K3v4/V9W2HseVEgDhp1jjW501FDA5s0M+z2
lMT0cnXFU8C18bUAK9B8+E+rrjO/UXP9DTCEfze831yQQ0U5+h/KlfjBA9H7i/K9
3oHKG80wAxDHrW3JQTObMe+ZRMIUGwV2wS7n4joRTcm2S6BE0J+KxvP29JXalawX
UbBzjceNcZ/M3w09SiveTeLLhOrmalHtM+HyX7mmLTE4bkQ1RvZqI2gg+IlV7tjP
pdPvUXJBvbU+Z+nND2Bvpd2r3RqrNRAGIe9aj8iRHZC1k7RSzr3d9aa/cX321CGb
GCpaef9lfgGT8ru3OqhvOb+jdhKzVQcMNnLP2KO1AC3ASyZUdWH7VoGzI2Ct+zIp
TynHL/W5Xf1xyYeJVAgGgc2M6U8tTYvMcyGKqPZRSXwiAC4dRDOIvARvdQQc9uxa
i5iYcimAF+KxYZYHHY+WlPfSf52UcesA6iRnx9ZgvUupbzh6Ft3oPvU4MT0nSNHl
z6OlUxUx2yWvd0lxCPzPHXAH0HbwjXdsusEDGyT+aJXcybFjtrZMAB1Tj8GQD3lY
hczgwEatBSlWcb0inlzNJqMwtWXrtUI1RcJnXVFxODqakVMhtMChvmAS0gxH5bI5
ywuoXXb594VMt+0vQ4ZkjBrLyLkHiXq6JEhT+d65R76HeGH6Jz85AD031UuX7wJf
kufolU9smCoHwQAl5odi1wh9gPZ7XKpBVp6ER/w+Kl6ycv0YqvXkAHGubq4VwhzQ
NJKnPeZbdSB3vGNObDiH1mAurd6WH239dLcUJbhfcxt7ROLRFYNuaZcIMywYjczP
eTRwXSiTaAjv8l0b4QNOAQXooCeTztUkLzFD6y8Dhw2OcHDuR6aqUsXCqgV+Fj3c
7FEEN5MC5PzJfbBRa8xP99JqpVQrw6FmHRKkJToKZYHv0dh8gcNOxyxEe5bI4JtB
yZpzQnGdWASn0Jfgxv9vrTICUZMFTA/82ksIsvBfwLdgSSYFE61/coDCNdb6+Huf
qn3qehGuAZ8qunBx2FFyVS7Hwa0AyIF09d5rBzC4hPt1XnQMjCRjO2/9T07s9QbE
AMvo6BOulGT+CEzqgvwXdnSmGh3fVJ2agmQlWdB1S4Er7P1UiWjdGGvtsAwmIRjo
MbsNY+j43IzvDQ8dn5VB2qJhK8TZhoVEgX4fJDFLEQrcAAe3KHyunbwEeTC3WAzk
wnUK9S4QFFuZoK7oGiLjm6SfnrSESx3hAL+dpuYn0woDM1NbFXgUUyWQQriDM01Q
Eyq6+9D1cwZ7opDGmsPM4tEIpcpgsvD0sw/8hO5UZLeRLam7LDZOX7ZP/UFSAJ79
+iC3boSljMguUYWb5I8cxX+I4p4q9WLAZm26zpaxbpTR+vJSxr3XEFbWDJSZ341h
naN43a+OPjyRo7Rkl0SmZw2ZHb3QC/f9B3z/MNOa02GMfJ8dR/2jpMNAPFyfVFxY
a3+a0WTKwpe/DlHWUP9pHhw1pMQ3o32Jy0Q5f6TKjZMmpHrOvpUm/36SyLg8FtUu
Sp9tbAXV2dZ1+OPuc8YJZiLCT9J0g6itMi/EY32Xy1nNoee3CfUOD621T12uNKXZ
MSIJJrVyWEuFSf3OfQBC+Ga9cTYKBwMP+jqH3Olw0HSLMmAzvw48mjKUtkbS3hpI
/P+2d6jdI2Bq0U64eDEPR61MS75KkjaP1iG583NjwVGBjZVsSFNPFQfmzKmgDHce
h6ZroQ+HXzffVHcJVKNeQx5qF8OOw+JIYtgOacmwJsMO5aVXGfOmksS6s55mwpi2
RqJxTu4QitKUgltJSOxTZ0irKalJjnmPdILyQNQy527tvIoEq7ESW486Ap1yq4xC
9RpzRtc851Jm+HDwV50phb5FiecrIwDj3s9A826gABS9FZDtdy4yOKIto4sTFG/m
ycGBEnDAEkVPn6SDiMeXlwckKIudP1q3sZ1EzEIUQEXCuM6mQy/0v2eQli3GzvrF
Ey5lmJq+wWp3tlz93OI6YjxvYdJ1zr/vPE07RRGBS7y6so6mZOJvI/kj1RXKgeK5
pBubOCpTJK59XMwfN35ZQcTuyHPxd4QD5Cqz//fJwgEPzlpT/Vw3XwT+eDN0X3l6
YOOX8GuFmgPln3U9I1VxguqX16PWDpvF7z5ZIahfFkXgElL4DVCoanNe9XWZ9d9X
mAvonTvwNoCZsWDQAe5uj6SSRH+Bg/fi1RFgwKpnVSmctgynKTBEvi1tXGOXgq+P
sM9DXHcFVlaKMlvZpJ9B4qqHIIXumonYtaM2GUbXDc3J0ELQXnmd6Y51bxZGneQD
wlHns1DUUwzBgSF8SuH/+GjjgpfQQexctdeo5w/jJZU=
`protect END_PROTECTED
