`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H4McArRjCFZjtsXxcFaUO047SbcMIZZ5vrT6jCfLpnKNDKiERjFLhyNgmUKbdyDD
ITgxzb4ZeickLM+1jeGiaLHxg+r4bymxsqLlPT58h+s1UjM0SHSHoEUQHm5GIef2
1mbSxqU18I9XuOBegROqQVb9ZPGWuOgSw7JdC0KgILQ41dyJrHbvL+41TXTUy/WA
lmpB5vbfizc0adDT+WwXxYugM5ERtsabYXdHeXzyFhHoYTrosymWssRpZ5ADMnnr
kNg6IukKQ8xGMBwTY081qt+kvrHVeHGBNmFLfFbmBILe2Wpi7wyj/ZAo7vbfOceH
QYxLgxpzkK2YElE+lzT20Dmle6RPlePommJ6ezBAsR6pKH/LDgLCUIEo0SJ1RaYw
peLHbDM+ZrTdg0F2ocd5plNCFsa6B3Ow3MKwlEaDnuTOOwUtKoJospBhHVcCW0oW
KMo28nF4iK2z8UkjGSVESDEmZEjRUm+4VsI6lqRQT75O6kZmR8lOqogZGJHIj3ge
pMhOOFDKKsGHhKl74jsJKXupxIQiMT807UwghMLou8arTNf6zLry6JhJZFpX4ASy
Qire0t0rLb79ZFJ+zLAjUIddaHXEUzyK/l5d/EkS5Efdfx6WxUyKqryl3hJK07WH
90WcrDuMce1zDfp4nwb0EVela67yF48AENVolG96/i+FutbfmyBYmSvGXT2Dgyf2
OF5t7v1ADFcutKUa7A22MrHdRFgp7Su30h9mEwowap3jSbTRikb1wNca3qARpMFp
`protect END_PROTECTED
