`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YPB3Tz39WqM/JSqiPkdoPfXpvYAQnXaGJW5aHBQ/wHT4tqvgT+73ruVY6ZOliD7V
Kxscr25gIH9CwkJCxkhOTfUkG7RByEHzbZBfJ9+K0Gyo2GtDZczUUej4afCh8lWP
c++Qq5i+DVKBaSn6QwPy9X2GHEDegBkP+dWar4k3PTxn2h0vX4ytPPW5yHkefyEd
8frk6T8DewrrRuo0vwl4aiAKLa4KwyBuNkx0VnoIYLQf6bN6mxJcW0wc+5bPzw/D
HoO/nK9dSZvKWWtgKSKIIta+F2nbo/hZSmFz4+Y0pXk4qPI/jXvuW+DY9wORGDIx
iftAFFPZ34aollNBwJBoM8TH9pI9ejIRitDt2G2eBEcC/iiLEwHIdNb40TBdi9lG
8ItAmbVbzbt1Ch68kxdXi7RbvIEqEOYDo340era5lQ4dKFRm5yUUGDidW06J62Vq
FhR+HlZp7pGwyQlowS6Ir/iqsHTLdvz1i043my3A5JXEpgZ5l/mIjVrFzujQDn43
D9nYjW3RkO6Ndm1zGJWJB54u5iEutR9NmHXABj66Z8V6g+qf2VLsPxWH1agHQL3K
cH1IJdWCPs20yIQGhBnOjnRJTmg2DntFCpo0bCKmMDytD6ORsKcmj4n7nCF/YZLN
Yia7fpe4CudwoS/RWlBNC0SNo/OcO5w2vMsoy1cmnduNhk0MGkwjLONsDNGr+13O
903ds5a4//o6fcDMJ8M3fc+JL1abLvWiCeZH9lq5uEnouCL+tS5KHfZtPny1yiHc
T4A+PUy9eMrxIgRnId2+XwfZ922AEg/QRMyw9N6WWb/yGGBWsK7Ggx1lxt4vBHlV
9BwhQP/JEtCouxrbWIhU5PFh30WT1T4I5l2KtlMabI/86XG8SKwZaqyge8GVYo3n
Pt/LycX/Eg9rokrfRv4hmiFUbhqwn0oWKorhLiwi86VqrsB33LcFz1u8qaqYkl2O
5twMmvAIdQbjHTN4xUnKl4s1YDmojJIp2sVPUwXZMYYum/koS3f8w9EX5SoPDu8P
qCySh9yVg6zzDGav/ReRcaK2E60W0eFd5YUGDYInfdbWu9O5y8bbhmv/RIQQOcXk
61VH/UzHnp7JgnmjUsHhbN6qChwbVHoQ+EtAD+adegK8rjQUc8WwlFH1/KJaXDLh
hkpgiC6RYIM5rvrikoKm0gvLJtfK8SqWfFLQ38jRE7SdOOZWHwQEJVM7oCRcUFvg
F4wNuMV8Ta83ltvf77IgOdMB5masvs6Inw4aKW3DnEXm4stBfULhmNBO4FOlfWl/
xZ8XHkjM2IrlBCXexGcKekyTHBzB/Djlk3mcK8pp+uqhCYpwFg0iBJXguS24Drgs
ZpF2Zok5bnonKp6OfdAxBu7+xTMu/HlqABgvIjFZCJkXsnil8vrvyvTEiTr5+0e0
dUy6rydtS7Y68pc7/5w46lI9m9G7buF8/1m/oYyTvxz3p7UCtoe4g5YjfyYfwUhe
//QmVZTGGSIXFvMyPI9YB8H2OLBYJ/X3wpYDQkFRlx3PfRAmJ9xJNWG6A5gwcsuV
inoNWobyLTu2KBZP6xyUQG+IoyLveUitmhfbqakVV0usLG62rhEIGbqE8+jZWr0V
TfJzQ0rvPBP+C2T3DBpW3/bjspZuVubPmiBG2Dy+hMmDST28XZz9+sUVG2KOAwQR
5Gc4LXq8l0EyjPXEIqNHbqz3t22gJjbkmbIT/YiG5xw1R72Pix71icj1WjOAP6oW
jHDESo7k8hfSfRnkRpsVMoo+tXDu2cW1T6VNSczEgeQzsZqhlVqKitE+GsaTv7y0
`protect END_PROTECTED
