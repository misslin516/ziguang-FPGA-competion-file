`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PyuzRMVh0q3rSRmLmxP2LMaM7tuQAosJG665dnHPqdU073oGlRxop2YTulOCdU3f
y1edt9GPMu56J0STH95uOrU+r/6o+oEPWF3RRZqlED8K3wImqwykM3P7OtOlStQd
EKmmsQtYSYkhlkB8a2L49ZDtnBT9jHWkHan+pEY3oC3T3qkRY81AlVjGehhTB6em
ZJFhaMbjPqcn/7pcwjQHa1oAeUtMocO+K1LfQcJrcL8kv1efGM2gqX+Z939thr1b
mxJqGzvIFZMLh9SM+aHdmwQ/bHfRF7QyklbyAd2kYUl9Sh46nZrQ9PjkE1bODe/j
mAxhqBKvTD/AqalR/qOd435e9qhswS+Aa30s61avbisGuNkbmDfqLgh/LxNZE0qj
KCek0JBZm3EpoohN/re5G8/Aw2uekLSir4z8QdoWIqZp5IcG+rm6aZZ9YQwnz3uB
WwJB0C5EJwNNRgYpUGV6Igqc1zehy7uboCbPmGSqOHozy52Zht/IXipUKwxJROa3
QRNo3g1yzyZCWI6GQVry3DJ1aokKFJJ00FQfXLF/rzgCrbWJdvldc/+U+B7UM9M2
oIap+SBlvzXHStorHo1wQ9pXhFUYGY2GlUie1APM1LKRJeHc0iTYX6G+zjVX1v49
bKiG+XaS6uvSc24mffU2RFx6laueGI7Hz03T+dsW2wYobwXhvWf3HFYk/6Q8NNrB
ny+vShAwPT8ODJs3/af8oGsQdPEjKGVQH8/tYF2kdct67dgU9dZUYN2y9AMWutdh
aJ+OmzxWoAeKiIY00eVxew==
`protect END_PROTECTED
