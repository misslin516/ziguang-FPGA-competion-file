`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hnBTTlgiUeBbdoQmnv/cSUIx7vJB65AhvwaYxKCCxySLaURk5Y8QrjE+/PylTyqr
bCgI2TzI1RGBbJbOaVaWoLbSPjX0vODUdj1+zwhE9PJLTuN2QdeLkR5fiex9rPNm
pV78uBrzoMqnTUDPlNxnLkPlZzD9eDQoh/M0uNNkRP9xNHBnWYTKUfJ8cDyz9Bi7
PwT11HJfaayYUYgiVrwQTKmSeeR6HoN8/cG6qIsNU5arFD8XnX7CZhjYn3yvhDxU
aeINHlvOV9gXvRnq42OLpt43SxqDh1LyGfzX2KGhiGk/WPAQL1FI+DyG1IGvJUVb
TgPBvokbbU+7CAZIbY+FpkwDMnhkM1jK2MXLISLe8m28OOkNDvcZkOy3NGcY6+sE
eQachs3PbRFf86imjBkgfIwtfFcABzKGJW7+n/6y1SjRySnRtX2KADZiGciS9lJv
4Mx46fOL+uUc55Tw7j7nlWZMgsqgk2JbAiZ9B2NvOjs1TVSLD37FG/YDMGh3qsRo
baDfuuF/Uv1JizYqiAFKJ5mdKcRo4F4NmEDO/Yj0X2vn3FCTPLNri0OBDtqjufh5
BRGS5RCiiAwHCWWlpo8CTV+ryNFS2khAs+N96nt29T1Ju+6tdeiGw4+5LDof4u2N
9h3XcmSEV82kkMS2xYk0jgP+q8VY67WF9cm5McRvXHx7Tf5wb6ClG+m48mjU9IKv
XdBR3TWy2DfQGdTbUsPR85x7+KiUe6qfdlRHJMXAmnj3qhlXxVzBKpHPvrjL+t0W
Ovk7SknpiAP56FwtFYc5pCSDx0VDroa2hDxJ6B/7Ut2Art8MWfZOGacWlfN4ciPW
siF6feNTJOh24iJsqdGo43PeXkhrkaQ96MX4nln2xfY3iDKmfCr5gf4UUW2b/56/
e+1iIfSSnOXa/TKCy460yB16pf4RAPzWagfWyTT0uVTZ09gVL0kK/8+xq278nYEQ
uQibpem9nc4cdwyP+ZhBcWNzQmQHgfgLTFuIg/e6jsGbx22HgyCvNsxk4fdq8qZC
wFIVd4JyEmau4YaeolKnL2KvN8mmodfuq2ZHAEc97U0iU4FfG5tlqpaR6scTXxKL
N8+zp1hH91CB/LuLwbUZ9MT+ykOhhV7Jpz99gUUp9V3ejimYKQL3ve8xH7OynHxM
aZo2ndvQ5KAvPFO41sM7u2c1QVYP/506nXbX+YxMVvPBfynygfDbVNw9E7ncBFPb
UBTUM0MXsLjXLktbAhQoT3YnBIF1nuZwhvccni0JU3BEd4AGlr+BOBb6b+XlHJtY
MLDHekQeDCOUtr/2F49INdHjSIlhgBEMHjGXlU6J/nxt1JFfsGVh8dC232l/dtpS
HWcxCZMd8cld6EOn0b26UW1IZ017e4wgS6PwUdMziG2qf+7pLGuYGG1pxOz8nh0d
8Yfo/M0Mvcu7GN5osPYC/PIuMmdhVWAhe9wDS6Pm05KNCTCUcVk4L8T8y+D35Lh3
rt7T1jYl0SWRqx0Rm/PPTOX7XXtD1vcrEXe2RDEaCKuBvP3hEMfK6Iu0QxS+YuSc
CPJreXW2uGdvzfp4t5hzrkH7M5NHPa+dcu9ngAnjArC/i0GH25n7MqwMo3vhLhfX
u9VQ9BTScV3NvCmab8NWzf3nufalBy9QJLvc5nLN1q+QhLAarcOkEaZzz3wHi8DV
2Kxz8g4JCM0zRmC3tSnveQ==
`protect END_PROTECTED
