`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMRoetdEro1al3iisobX2K4Ex8R7K7mKHE7x51Z0nuXU+Ym8HTK/IC7ed5EY7sss
io/Xw0cFeVdYrl96i8mjUOntXPd4NBgDmRUrR3GYfKOlSsTRQnzcyYWj0jZxOopk
DgSZjlyy6hO/leKgO37mOIewDLi5MXOhbD65jT5Bm3xKeg6q2EX/h4q3RhT7+6QJ
ceBMd4N4QM6NE+5aAj8kiKXJPank+6miMk2XvX2DcIXpQpdtvBNyztbxkJHm9fR2
JzEmeJfHyRoYEqqQoYjl9HkqeloiZpBSldccni5M+370Oz2N7cVL2uaLsZO1RQa0
PCvzHNOqPMB1/wAIvmAibmb5wdlwAnJVIECzIKhc3HLKNjRm1E1Mnv5XTuT4bfO1
LFeXKflpfyCb3lIGjGv4HcfGkI2ZOgZvBkG4pEsmt8heQDExS67wuH/+QiGkXhjw
pG5A4Rn/1kG2CU/WglhpUZEDPy+1YU8ALK5frTbjRhGA98H+vGFceIblAdQbYm5N
2RoIwA4DPWVbCehsPNDHoJVS4xxvbxjZbxq3LiGvyqK1aGXviK2MqS9yqE0hPFIX
aTt9MkAkAF05f01AHYu0GOxTPeAFbWdvnPp0YTz6Qy4cZqCcni+HVwD/x0uvkazA
ET0Bkp1oQjLprtJB0O7RyCOmi7oQ416bpff+7pMeN7DapB22A/BrhaGucaJFVwOs
dIwIgh+9+TVz+twwH17+rwRWf6VVbJ4CuDOG47xGfj//wCirjzuPkOpEyuR2DGsc
0l7visOfr77AuLC4Mxo4peeCaJM9jc+o9MxxM5LlDhGc0hEbi9G5OgLTRMfZ6aJ9
xiGVW1NSTCZ+uEUNunkzC0HA7ltAn+Qrwsa4A/vDDM2FmbmRK+ggpsB52rXg/eFT
mwAmgd282BgqE/nAxBVuBH6yjnqQmkwz0fei2ZD0bp85AVkYP+0Uh3gBL+ICD/+h
mp7MrMlBCsdiGIcm/Txwnc7iqxqEvU/wF9go60w8+ZeTff03g5MHuhv7feH77kTO
yokvgj0gny1RqoQCyXAJ6PHwZDjYkry9R+1OLY3W9WQft8bbvJJlkQyiCxtChpqw
dU28YRxtjOvNTJHx9wiSpYynmcYY57llw9mpzcsbM+mYpvA+oOrLzdKX4ws9BlcT
bjvgEP4JDUMe+jXM4yi52J75Buf3g5dg1JXlxaha6elStzxhU6wfF+e2j61kars8
TBKlRrQnPIh26IKvBhJM0UyBl0z71hL3rFIW+jIcEWKiQ9JoYaoFber6Fg7YMWXj
mwRfq2GBLh2qGRUdclbZXYI1VQ+6jRKWonpT5R6EHHvotnnfc8++p3b1x5av1Wfu
WOXw15wIEXxK0Cy8AuvW4Jsw+BM6lrYcr0Udo4DkyeYyPlyBwQRwif+d6tJqZx29
KVd9Q90VXn/y25p8dDncvr3lz0nhRf6sNLUajPXL+GKdJty/CJfKnyBo+nfdjDRx
+ItPiLT6BWfZTaKYD+aPv3e9SXWZbqdikw+W3PNCBOz3tNA7GRRxd1QQsOuIbrLS
D4BjSK8J+jzgx2unvnGW2KVM0xT8Me4y5Jg7OaZQqjbNEf7LTeDIod8RNowybLQ+
+cO/swaQLG6Je0IL2c+58PTOkhhr42l0/IJgiBpBO2aq+o0gksQldGi5/AFZcxcb
GeMhsnYcOSgUJjCgRVqEJ9R0hbItlKoVrY9jRUiU4nV5Q36tiwVBBKOMVre4UEL2
z6fj1kI33QT3h3B/8MBW8Qv8EiBXY9/DvedXBwhKKgsVnleiidZK3Dokgrq+Gf+D
Dh7vBXn+c9s6LsWfh+Erc207a3DF7M05toyplKtvWPGmYI6LWtIpcykO0dPP0pj3
fC1DRci58bl3aBct57rSc3UGaxgC4Cxiq3PZvHwj0hi34GmEhbrIXSSZJ1NtoYDv
ePAp7B+k8uZXQv13B7NHjgyp4GuvhZ+j/tSwP1hILHRdi8xGwI5g2/THKuRGReHn
bzrVbkXVqTlHyFGSW7u9lr24fKZafAnG3z7iFIvjRLXZi8OqtZqOFN2d6glr0Kda
Qf4c0SHWyD61P42QVKqhutGnI4aiT/98CwgNCxzLRrtk3RwwR3p0uvbfZXzV2YT7
Ou2qyU9RgjRhvUDAQQcBEgFVxJRCynPNOca13A3VYf2bTFF9dTqHxiRjTzZ5NBuO
xeJ7TWDr683FUsLkjYxqn/6OLPrEoW2HfxoCXVd07VL9iWzUVqdN7ycMl4lHEG8x
vZT0+L7W5v0Bj297KRAx4R6n3/bpV2uLHwd9Oyv1qwpIZBIDsPEcMfbRvjE4YZWB
y64kMxuWe7i+pw26/EfPWjnztmL1rsMmljweC91jtI1AmueuYodxW35LA+ikS/kH
QX2y6XgQi5w0yMLMAohHDN24ACGafT8KY/rfOLWsuj3tdra9AcdXdUI4KGHja7Ac
LolpZn2JZJITcMhHffyyiN511NcSZSv3pewMODjkqFCcTV/lP+WIueYEt6Oo4NHz
xXm+mpeNifi23uSc2Yo7od20MKvJGl5zpuHV9CWYJVYDzrLM10KooLLASAMxhN8U
qfH2kD8rH4ZGV/+65ikJkzJ6XQGXcfp/eljYzN2w0fvCs1Wl4wZl7sSMHr4V1dcD
i71ry7XTnSoGBCCcw6TLV9hVWe5WY6YjzKNWHdmQ5R9CIfgeRZ3xo1Qkp1tl4JhV
32ESD+Cggebd0CEUn8rDaA1HnU6sFN3Wd3QaUJ65jjKsgcBWny8ppUK7Q8pUa35T
prEw3l9xn0lNnK0tDTQ0t5ILp7O+2lJtF1p8Hnad8lhtueHebNH7+N69FnvMZp5e
4359XIb23hugKOLJWrcTqWgbk6GQwWEAHqf2x9nIGbtFNV2HY6EagVS2UrAOStp0
ieX8qH6zfZPYpdz8a9kr3HzTrY3hurS3EPnGsl1SzSEZxuoNirJVyBzeEliH14Hx
r5M9Es0mFXLKORijtzlgCeBAfjFolgw9NltTXmf12Lc54NPMPDSQp4MpYZ/50jtA
Yropa1s2MdG+h+jAG9pnzaxohOJ/5mvcNsUFhynWcH1xkPlT4hqT3GmEJCz+KmAV
QUghH18bgtEQphP4AMNGGH5L8XWVV5XewKJs7dh1w/72mSgTp00i6l/EaXvQa1Sl
3T19ezHh2ifa7QZsdlvdDaNJ16uq37lGC6/mAfwGgmvfe4c0mDHhRVmoZpove80w
646rhPMv7Uc749yQXD+3sAzctfQfaqM3klXzbXvKyx+OadvUrjnKLVeVJyMzQTto
EexCJRhkGTtnAMXFL/qI1ZQIx82B8kyQQOeWzyjLURFKvSUOntthh+eAR95Vcsat
W6T7WH5c1ZzaEuyALXJGBC6I0N0232t7ivmKp9XJQwd0k1Lg6Zg41RwtBWDl4eGc
Jp5Li4bKGOgDCRKdpCrwnVSP0UzZyiGYYKIYhDy4hob2Z0fRe/a+97HJDPEqZZEC
/yIWFQgu/CtLHqfLNPirHvRfjAkcloOZzS25GH/kOtGadK2dtyd0U++99Cn2ymjB
SbcqpnjwVZBZic+Xkt6arocOsr4H/ITztdJf9dcBLbiRVmSN4pf5G3+rYEyzQfFD
5YFSnpDKO1Kdn5hIjKeC9RP+eusIHLUU5H5kH2wThzkQRYok/lSEXK7TgJ9NhJ9H
7oJXE2ZvQuvgCGU+vaohQgyDKOUuTJo/LSxRUx+ft4gT8nA0nc1Y4dI4IE0H+1Ax
PipxaoaEmlF+SaEYRbAo/PDJoeyFWN5LJnJigD6vQLkziIQ6XJNNYFSoIyeKU5eq
jY6UyjWFzfBPnTZHdeYS2xJyM8KfzZz3MADkVbpsq1i7bRS7JaHiWjXEyGKRIrkR
0YDjxcmljJ/haAez/CXscCCT+g4S+wbJBRnBcu3bXeY8MXERQ1HI89Oys+9OlAsJ
xf1SGcnyAFpYBx5qWnbjLvhlsPhp6c2OHnqg18hP1qybJGpRtM2OkBPeKRvUmTA/
iwIFFh/kT1nHNLCvOEdoqP9s30QY89LQ1Em4B4F0SG4JOh2RakZi6hFAcX0dRnha
MeU6gi1/Gkm7U0+prBrMDc1aFW/SKsF03qAMKCCWHGbuMw2/evj6OJ24l1I6W9c4
6uIBqpuTyf5/szirTN23HC5QKZPswdYFhthLMaICUsQMeNpYt6nHBwL1Gxtwg4Eg
GD0Ye+FAORjEvEra12xwA2Zmh47ox1Ek5epwXQBsMjjzF5vcEAn1e2yN8hFbhQNH
WDjxyEGbbpygjaVy0QcuJpjJ5644Z7NfDZMO2v5xirxFB8hKlgqXDdIN9TCVr3hC
oVPQpI+p0MmEQ9WUbf4LowG7VN7bGDNajZooPd4wH22k3e6LX/CofAazj0CLpViL
Myc4ltI/DY1koKTF2YsxOTVJkALnxetnElQMD3ck+pdSM0W8UGNCdUwKp65gykiR
rJl5Sd4jvC8Ac/KjPAQXmTs+MpcgO/s5NT+kUZUhi9OgMYXt80pATCvksL8T6XLu
tdIBVBmMUbIoyatK8LiECY/FdUkGMxwYLT2HbU9VCwnQQnLCT+suumj1/9twvHP0
OAGz0fJQduuxXg4p3tSTEZTs5OBJqZXzfaGH5MivnRelj4/YavGBpKClh+ujpf+q
SuODpCuMvtMtpFrqMUb4Ai8yRYYDq4D0jdTvTrtfSR6AtJznb4JmzjpZy0Tf7QUB
tBwha5wj7/xN3ZWTc6EkxnqmDYKbHLHSNH0eP31BcNRHvmRywEl+FNs6TBuf0gt8
KGQgTC5dc+qog6EkQ1sSlvtSVCLxIVBLJSOvwJWq4to63iR+vNuSvMML0RIu0ex4
gQyUKTSxKCOx/f4uUQaVtsOj9ShMM8lXHxbiz46EI5bKZ4rd4sRpcc3SpeBV3QwH
Mr2YPchTfosrbyScbrflQ0DVQnsDVH+DulpX0zEftg+5yiHh+Eci9SxskscmGtLF
xQjqkxCMu3KuLCjMVh1SZPS+Jy7WDOPXH/VehBQhYK69stoblak//+YlPf3HM1FB
x2VQFuBqTjbKBfBubdHG1SlyJ9GDiu5vCXbSXMBzbcx9ZxhpaCGsGBLAf3ZI5iTS
hUHPJdtciAa4ODc1/oqiDE3DI5IdAY1kyYUd0E503MYJ2ZIIhuSE4mfhZS71oXuO
iSTX32MWbfZ+kjKRx2PwZwpwLu8ODkZW8wTTr69H6iOn16ItW9O+J3rm+rnTfiOQ
WHKkm6tijkUfRivC/PuF1rbAfK4pBiAjhGoH4LXjzmPnJ/moMaVEhu5gZJSuHdRx
YPfTUAjGF3cVPXKnYKtor7VTTWs6bR4lebVThQdtFHs=
`protect END_PROTECTED
