`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MjAfwCJ61CT0kaqZxmGVOHS1R3/Ix+MmUccg/aulrTcjv9LlMsowk0sFcy7atwxD
lK3NC4E8AQnQINyr4liLrcDNtyA+LQaPwU+VPQj/yaG6IxITQQSLJbXnOtKNDe/U
clx7G9zGb76VSb1abCBJBjMN37e5YsKdLCHaoobuRE/2HFgzzD4LciRtFDnHRlqG
qhOv8yZTiexF2VRj4thBQcF2gLvv/6fX2YOnG/yAQa/ABWHQE8yAGQpdquOrJP5d
Oc8YbQF2AFqO20AJlrxIoiIPcPAJJNi4/s/QAIiN8y9NmKEVaIt0dxOvUhJq0JAx
msETPYPTPSlsHfMySoiC/iLVRTZzlJmzNfoKo3i4/cl4h5ngAX2itjzmv1zliCF+
LyAp1EAnZXqm+bJq55zL+gbDwZtjnxX+7pmpGzv+zlJGyyPyAkPbWzdBNWQtOEfZ
txLax7OChPZlRdx14ikGdmw/udrnMUfAc+yu4gimX6MZhsIMnGNodbiFD04wEtLg
3hP3OrtPgZHrqS5NboJc5DdQmzlZdDDWRtbj+u0aK82Rjhf4sdrgX5vojPTT59zm
uk4ttmMUp10jKHdpnry7V+ER1RsNsr1LghhWQjFQpAQbbps1z4ABXps118ITVc6f
EAq2Yak1+OKEWGeg2UBbpjSmY2BeXjDQ9ALXXiESbemGXVLeVohepLbGoVQ3q6Lc
3X+QVGwzrGbH2FkYp8PpkFJLae9485WIa37TnZJWapYPdZNUFVpiQ7dUfgIbf/nZ
KYkoKV+GhbktY65wrWX88Rh05hqiGDzQ+t+0RjeJnLuQQEl/w77AJqJOWEgrMEEH
7JzsoUzWmo7jJW4eCt1gEtPBehthbC+HQ4Rh2NPsLKHaVBKNZ7XAWX1n68gsayau
xgrN1UXuyBIFVIrlHtG+anbQnooD7DcFpoSaPlVhJ8lzWZs+V6+hGFE6R0EqE/A8
K1aAs8yr2GXZcCc7StYbj1YUdS69gR/RZ0G23j/1kVofpQGxSmjknuIZABlFYsQ7
xETbY4p228X2LNJXk+kZtjS9iVvyvjrFtBwM1uO3u5yk9+It4Fas5cSAU36gBxq/
yMgvdmhDhJAJ4vVZN57xqfCEo3IAGxkv85VNHBjt7YU0ay39XwJQd3hHEpHlUCcb
LIkeO37hUiI47MYWx2DBlfsbYt+EyEvDzvkrtgPyk6Sxvy1ZV34cScLgTLOkP9aJ
BnY6pul8NIF32N91FEw+SUKbJ39yLg3+7tknPEtBQI9HG9FAOUE/3l7q2SqrBbs7
6IrHh9lSh0iw4hyzvfqjL1YRVCbmCtm3NsZdXyhgcVA=
`protect END_PROTECTED
