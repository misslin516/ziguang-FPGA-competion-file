//created date:2024/05/13


//*************************1920*1080@60Hz*148.5MHz**********************************************
// parameter V_TOTAL = 12'd1125;
// parameter V_FP = 12'd4;
// parameter V_BP = 12'd36;
// parameter V_SYNC = 12'd5;
// parameter V_ACT = 12'd1080;
// parameter H_TOTAL = 12'd2200;

// parameter H_FP = 12'd88;
// parameter H_BP = 12'd148;
// parameter H_SYNC = 12'd44;
// parameter H_ACT = 12'd1920;
// parameter HV_OFFSET = 12'd0;

// //*************************1280*720@60Hz*74.25MHz**********************************************
// parameter V_TOTAL = 10'd750;
// parameter V_FP = 10'd5;
// parameter V_BP = 10'd20;
// parameter V_SYNC = 10'd5;
// parameter V_ACT = 10'd720;

// parameter H_TOTAL = 11'd1650;
// parameter H_FP = 11'd110;
// parameter H_BP = 11'd220;
// parameter H_SYNC = 11'd40;
// parameter H_ACT = 11'd1280;
// parameter HV_OFFSET = 11'd0;

//*************************640*480@60Hz* 25.175MHz*********************************************

parameter V_TOTAL = 10'd525;
parameter V_FP = 10'd11;
parameter V_BP = 10'd32;
parameter V_SYNC = 10'd2;
parameter V_ACT = 10'd480;

parameter H_TOTAL = 10'd800;
parameter H_FP = 10'd16;
parameter H_BP = 10'd48;
parameter H_SYNC = 10'd96;
parameter H_ACT = 10'd640;
parameter HV_OFFSET = 10'd0;


// //*************************640*480@85Hz* 36MHz*********************************************

// parameter V_TOTAL = 10'd509;
// parameter V_FP = 10'd1;
// parameter V_BP = 10'd25;
// parameter V_SYNC = 10'd3;
// parameter V_ACT = 10'd480;

// parameter H_TOTAL = 10'd832;
// parameter H_FP = 10'd56;
// parameter H_BP = 10'd80;
// parameter H_SYNC = 10'd56;
// parameter H_ACT = 10'd640;
// parameter HV_OFFSET = 10'd0;







