`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HHmxGp5Z8cTNHi0bXO4Fflf9oL+wZX8RWgi0z+MpHQoTZ6S3Y6Lmf4hVzlKkAn6H
5azRnJG02Znqe/LzTit60mdLvmczm+9yJjPFPoXk8uHOAzH7oQGEsqcb2Hc6TrWG
RawKYVI+pU8Im8esLLxeCWSTujxCRPTrkz9pbbUtM0JH2zZV3Ygy2igcQ3D3oH3y
F2Bp9FDZU1syRz1PU4WJUr4F1K/qnp3N4e1w0JeLFxTqySoyD6IYLL3d5p4lBnxd
bQWaMBl2XYIOjFLU5/tTQo8qmLrjZjCqYGR586WV03UTHbvf4aVs763GNbJ6y4Du
8ySCD5K0unKg5DFwo3BeBA2nmTvgmaVFudkKz/4yKejT8pv63FFLFfgXYFz/CumM
Nj1/sMqsIU81GPdzTeC8Yr0QmJDRRXQO5/1ilzZ9IoPdKAkJHZ0gp8v0EScPtQUf
s8sBN7NSqZpemSoy7dNveoQV8/EJoQ5cgZwyIzvhyGlrJJccSZJzUxzXfyGeSY8Z
gNqI4NCiEIr/W3cx8LfyLg9cW5Ts1IeLegGIRJybBolveOvJsRg5w+7RxQq63d0W
ByYRMo/asofUy63vXmzWgmkAoP8a8wA0KlFMPPMrBKdaX1A1JfLSYSYcknmePWVs
K35Bdbu2AvdW3WfrnDKPS+MbinbLmmsS52kXGmh5vcZp8ecJsYuDDdoIYfdw16hu
sW9Fu97w7Ur0jzN2TRs+r9gJf8h7xRiIMBrwfOxIlTPJoBpWXXLnhkubKQQnPZNM
FXbbaZ92kwAu2rLLApLsKauXOuM6LNvw7wybi/1qMUdHOEBZlNoSGup69zfQHoAS
a3FBmApCPTH3djEZPCPN+YuVUQ6IeB/1T9jSQYKPu5b37VUZK8bvlIQPNYKGW6zk
gVILnmQPJLrIo2oZnEEVb67RYQCvXTkfB8H1xRNSmjsyhplXYPJRzluTjt4g7RI/
YqCZeQrI3pIJXrYp7cZg+sK8GIfmCf0c/ORAz1pg5SVc+k8zE/S1Tbrmro3MAqN4
azaqoVc9qKW4CqzNcwUrTdKRFFbRURpYDSj1WPmuKWYe9mgmZ680IqnavzvgLNZn
VeWzFaQ6tHVaWX2PheWCSRZ6ic7SBHDc205pzcHiZPOz/YFqNS/iHOMGluCq2uEU
Bx9s/eJBUwAplEofwUaP1Q==
`protect END_PROTECTED
