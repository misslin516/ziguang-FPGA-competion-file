`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9iRrll5V6cpEghQP7Yv2rLoVkPIhygA2PZnxQpxI6ndRLPuStsZHfyMRw/a1Gqm
0bBKdfLm9kh5qFCxQFlMQwLDeadWrAvRprp8DlqAdWuFT4I4Hyd1Wsj0tgjlzcvB
yvsR5i0i1jOBbYlwsBde53Ta/TBx9efNE5WA9s3ZCTksj9cYT1LJ4zciHsj/0T9S
y2w1WXJH7pdbZAqi6xlZIkp3n70Ffeko6Y4bIn3WFeAOWiK2RnxiCEHQDWVdRHws
uGypPZPlKvNOy1ZjQ8wsD0WEaJeEOfZnU+4DFN6MBkwdcZ4kPOGtLRS2YhkDPUe6
4un7UZEKwyIrXw37t8woLykaG5B5W59CEQ7ob196bbem8ubva9tb4XSD4jDj7ySV
/THSf3g2CpB9Ow7XWb70FSmDgOvWDsNQ6gc7VN3rcUJqvpH97vsG8Nayz4WUDWf6
tfyvx4VYzYLT5kYeS/IoSM32ixgz7Kz3zWC1WSiqBbz4s+GPg8dvyXTcNh5m3uiY
ZwohNwyPJAfRtvvgFrPkDv8ThFFf8mAa7EdiZSvuIk/fxAxEXPCPEyrpHAiXmgat
CAqYh7If6Ug58Xk17p/KqAmIksMzLS3be8i8vJBcBTgcd6VKry1qYEgxf5ibcmZA
xN6JQX9/JdzRfE6Uv90Uqe4srdLZilyE62W388mqeS9I71Cz8v90zVNXGfATrbDu
m3GxImWa0a9gHPmB+v4BYJ2avi1gl/xHoN7Nuh9GL2AgBKqZI4ph5tWAg3la7dob
VyuuFvi2CwneZcpchleNHAEbLToWt7DYLdBkEPInvm/3j9XlNUKnhQDU2/d5sSSt
j4tjHXwmO54QKFKmw0oTJtuQJ/iO1GWBcWnEz1ugB8V7sw4//YVERYxw0v98C82w
uZzjF7YP2flUY7m7owhp6Qdw2R0rj2XEBeBDb/mwlqYZYAQV9hqibWz+sZ2GKG5C
03RkfGVMhiyi00F6NiBq/BPa3f5pgOzlWNmOXRqulJARL7DllHzjyW4M4td2QGQ0
0asEuigkenfF0XB9pleJu+uXMYsaf9pkE8Ny0WyJI9LYya9PbfChP89Jx/0FK+K1
bg45dXDIrbIV3Bj1RD6eCFpSv5p6yyF97Y268KQ72aejAkoisKChsxEGgNtOrQHe
c9UPOn4C+x2udLfEXj8d5ItvLjnNj9Y2KIubAVhfczSw3TWYruhbcvwdZy8gUFyF
/hhMsQZJzbnXsuMQJiL/b3lyxlxFvlYeGbimF7L8IKPUrh/qnRXttMil5IbsEeFK
nlcOXEMGuiRBrUGn+glRnm2MGjLLPZet8wiqORfVXYEHW9OnOBzvSqF1U4vvjMFd
kCQTwlXPpQ860/MVjQ4+uo/PbcVC3b/8g11aLpH+6owXJ+wOau1J3BszcDsCBppY
Vssu46dUEFCKx1Slrzm2wvtidTxi2eZSGSGFzQsqIlORu7VIDehkayVrpD0OOril
gPhItBm1HhSD+plx12MMN0ei0wIQ77rMnzmZohPGBwSN6HPFi9LOc5PU+e08OdNE
oPXLZIcdLNJHfyP5/EmwEk1UJ3ybHaU4gwH3+4e1AHT4WsQIN1cx6a21pokkj1Gw
nan9rpv8p1RrgbAiIrtHC67wXPheUzVbyk8QESoSFXB9p68Uz7Nmk2uVZM5DSabF
HVHfP77IuyHDAlWchV8mITcg6EskohWhkMmOR1KH9sVWc4GbBgHuTsBk6ehV5PoX
020NhpfuG5ppv5ktmpzH738rey0wurljXxB059/dE4Nmn/JL1ANUo6KySBP3SCWa
ph9nwCRHhkC7J/+nUcsnwTAzOufyEM1n2Qlz7CynXShg5899ZPL++QGT2uBwLwwv
WE2jfEutUpHCC9m7p+4tSwCFoa0O+kmIdT/sCXUuZOujgG2et2vF7kmyrqMZp7cT
dkqeMTTw63Iit/rXUXpbrtTejUTh+bhtx8wbES3uwAJRYbtRDJis56KZ8PRGhl5/
0Cfpn8tRpvJQsjS5Z5wjuGp+lshgzeUWuBwJsfTmei7qxoILZ+AmPjsS8QAfJT70
5PRP0svvhNsTs630KG7eRscad//xuFdx35IEA2bDqEWR/BFt9ZbLgrDHg6DuOUJA
5YrIxhnEckDpBypPViS5aVEmzYj1vyGbzbnSCnoyqvo7W0biNaXiVwIUZ+f2vZ8G
3GnlFKuyUVZ+618QHdvsJ9wsbZphLQIyD77AfFWd0QFM2knV+zKOqXQOdaPBS1B3
aGNPWIXyQNu5lsWdHQpJ/GpzESIE5txgvrRPrTx3L5JZ/2Hl2q9OOChYnqBW619Y
ub5/jShCOsGfG4G2frRQe6SUTAZWxRByxDT4TULppRydK/gnp6Ch9ZWq6p9w+qmk
EygxbhRSNdsv2fNsexzGYqnZ1UhKachA3YeEe4d+t8SZmdT9kfIlOPKw3BmdfaGX
IKvsCjSeOCB4qHfsV8b5KFaPI+/6KxoHnDI8KqTVdZPYjOjYvU4BjIiLDv+3uRqe
xboI/MCczKyJgGEcmRJdUdRaoA97HbmJ/ymEyvFhxzycmVJjEz86gWqAz8ROvqqv
gpyN8IIWvEGxATRXoF+5pP4ssatWoXA70BnKuEU9rZr97wjkNAD920QityGyzQV+
rLgczbcQTsQ2EMJ6qbgDEPin49Fl4RqV900JyXQmysNz6XE2odg5C7ETwxaajoO6
SHRTZxslIgNNOumPAXqJzay/W+11ukLwq5tDbj14Ykvnr5qUPTQ4GFFR0aQTBnMu
vDNFO2ksnLZnymiCvF35sJGKT3ejpPzPTizb4skvCwE773DIVikU5ehv+WfFAPiL
6QAs01mtD604JTPkIA5ug1uSGVIZy4Hl0+LnsBp4GXmHejZCms2SIvrLUmn0zShT
oNFJ1Gtcr7Jwc9MJbVf1F28vJWcuJvx+snPpee2NQglpLLgebI8g2q6G32H3keLJ
kefCWYt1wY/lun6VCUL2hsGHm2Abbg1zoTnOk/KRY/YzkP/ed4c1nOcJu5SbYIUB
ECcfuDC4Z+uYYmuuvfhNFejCNS3pxK8bU0jSvx2TUWCUldojz6JEaWONWPa43NiL
hDXvWEFThHwSBQzBmKmkbtrrl+tInx6K9gVWB13lHQ2EW/wobNekFVQjL+T0rwgV
61oswBUSC8jHquGznmlPNaYjUsHJYbdqfaKwcVbFE7B/g5y0el2y1573PvxaH4vz
Fv/V7liajpmXU5szS8js5qAOrwek5ojk4wDXsCfRd5SJvmKJSnf1vXmyJj+iwZ7T
FGCbtvPIsuCyg48MbUsXKp4k+ls1+l996iDBNvME7RAveu8TYyTjT+ZToOiG9lkC
jeUDsQK8W4fvKjgckNgoxRrTAwu8yPw0Itp9g2vWcK4RPiStwzw7G671lX5ykDTu
cDu+b7TY2Fli5W8eIxJ+9UZtMF8IT6e+Hsc5OURlrRIdyQg1/x2CSsGTWVx8pfZ7
yJzjLt8GntZJ1sHmD6HKHszfgX7I2hAAFCge7wuG0om80boEGCTLeZrZQvrc01Bs
76b3ST6u6v6HOkXWtr/jmaTB4n4bvgTAzP7P3ZFJmctsApcCppZxr0dbFYFtaq16
n/ha3PyrlHv5GBQeJhYP6TRYy1l1Zi0vuYjRuH/RWqgIkPAYsfoXsrFMubJzvvv+
G0Wy8yHDO0L983VN/r8zPSQx1KYPQY+ZeWCq1avOZlcECpluo3jdBN07nXpvT/1Z
41eJTK5NK/dj3A78Zr/UZubI7awbSHu3zHvtVRiwu//fzXb6qGNHrYRAV/dJDHMy
8ECcKqPlEwhPOjk3G3KCjm1qyUFzxgS9rMD0RvR3cO7btAz+GC+MipMON2SaLLf3
Hh+iTiNF1mTqpRkohEdRldFzz+HLcMI3w17kPdvZjIk2+R9tvYwBPQAJizxjwhBv
r7yNkvPYtERuXAscPiIKGshrg2H9iIPnK2pTh9FYxSExN2Tce4S/ravBIcF2iUPa
ImFL1A/b7ZLENijq3TZoS24SOyhch3Ck3ONlTxPxXb874vqoab2h/GTJyHncQpvz
jklugOraa+c5FoecqikNGUDn+EMOUS16Xs6gm9YmpsXCufXindfYvISJhvrdm5Zc
zwUYzlzVpW2GGCFY8uSVjYbRM1qiLaTQVjVpXA/wuLONV7CqWYdsn2qT6q0TEES2
xxAFtCl65SntTU7LLJdF8H+xAeB/DtrTeDxsWWkcJRKISzCTIi/aWkJhINPNt0Bl
uZj1crO58NG9+A7Fu1D3rUlKdiAwKZ9a1IllEGHK8qEsXMH6jJdZwAF411VmT0uX
XK9ntVkzDNfnlqH4e9bUEBzClFE+OCcTo4UVrFEcf8CxvOXB+Q1VPl0cYyOrWL1B
89Og0f1zviy+4bLsgRDg4jBTi7xUlD+uN+hnvhDciqjkK06xAzTN3XWc0d161iUb
1WIf4yH1GJzE58w0v6jc6q6sGkMfBGQI/kSFQtVSO/r7MoVQoHOwdIdXSxgfveNP
40BhDl27qcEcQDk46sfGpwiiQABd0mC3fJsabk+/m8dfJcYqa60RL/T+Lv0qqPTm
QXWnS8Ayino2eoCptj7FrksNH9kdYXncFKu2VrZdnav1QF+IZpzrBun5q77YnzmP
H3/d3LJ22e65oH04JCaOrqWEmPW9kEz0TOKQRDEjRYgQPLxNWcyPGFYd+llOqSMm
QnpHMWmLIkSgxTZkhHjcbGkX0RCb2awIjYPK0B7Jm/dY2JwABWOUXGJT5jf3Qpcm
bYvEgvf6cxbFSVNXaXeqqNjJoaXHXcMN92o/iABoIeTecH2eICn9sDVipwFaNKy8
99a+bNLdryh37+Kqik8esnAiWxN9tNETXCs0c4mw9rz7Tj63wtZged8szyRA2BBi
8PYI9gsXjchZ8miAn/acnyNZJ2l5zlRvbaFXKsgG4yfjs3ygVgieSOCywmwaT8qZ
Ty9uxl8x6+meGA2QnMFdDy23Y8+spKWQkfL/a6noy59fiSJ6xVgeB5/MmMx6PV4N
O19iLUMy5VPPyOhNFQdOV5UHphudBq+805iZ/xuMaEWVzCxfby5GB4sxZ0J8vVtW
8A7VYSjcdEb2naNPpLJVBgnYDMd/GmP1XHYGQZSOaHuo8Y53+NACaXErr+CBOEJ1
cGS97lciXhJojOkKXDgX9yA6U1+wu8gmgbDIXoNGbVXF5BUIAFj9frblTE32aNEp
OuwJK1+XsITWH8DlLO7e0tLX5iE5aSb/MaAOhr4pW/9XcSR63QmH5a852f2Ah+gk
L7ePtAiCpfp//26gT9fXqLuQSlX7zEGL9lt+NsRlAFznpbuw99uduOWEQbKeoj4W
WLiaxFHReEbEKBHsFduVL4R0oIaEaQOaU5apvitQauIFRcll4/MYKQenFri76wvt
TWt/rNoLV/l6OIJCbVXnNPMYzTl+SxbLoH9aEHQCIM785UzoMHj5zet/+TxGyo2Y
JZYMEWnvvAbRAdH4nMflqsgSL96t4xtnvuXFydUY6sMxbX4432JxQ95iK480gTbR
B8My/HYxUbSUTADnUgXiAYfhwiclDNd6nmZ/nBiEqUpZwG5m2+IAJsuBJ6IeOWlB
Xask/KsHropPdmyx3o618hZzMdXEc2jgCHZRepq9I8me4jb8BsPY9oZZRg/NGbRH
VzjfHZlaJnjK+wfCNdBbHdg3KXgZbXyQRUtV5vH1EA691FO1MkaStyBiZCI4dA4A
C9QeBUmbQ+JwkEwXbn/EQYo4CATNBxZr0I/aFhFSxRaVUuHoeFvNG2gSZMLXsLz2
AQe8lyVoWAI9tHT9T5Xd5+c3qHlLGGUn5XD0s9tS2wiIsCsXlHgcR7VdNieQZzbr
2WztqzwhNXHSgfBdPFQ93mY4Idorm9P/OX6xCjlO4ACOfZd+7+ih3wGCbwczFPEs
y2KzLZ3hXPgvU6afmRoCpcXGW+dWWXk1CNsXLqCOYXc6uQU1avx+lzRSObZy0vdy
p5/gfYl19oq0wKIth9yfEhV754vtQHOkAa+or4olS0NM6E9EHsUPzn41Np+S0+vd
GGsw8qFEDNgdQD80GwWX7Ue52ew4IQd0zCZavJa7+AwFRRRTK9nOJof+fb9UGZ1Y
ZBPo0cBUjo/+V8QdrHenkciRBTJgGhhgwFyPxjdNkt9LtGlsk0u5Co6osNCQWYox
+bmDds+eDn/UoTldpvbiBDwAsY3XDJFK/Al7P19GaRag/y40CS3bENc0zwbUkmGY
a3dekAk0xiJbykMmvDJQHOBcHuCf6MKLdh/U1QPqiXmHFSMVhxdvwb41Cgn8zIih
RzQpVOa3GdcSeQS17NFO8sKlDXfKMd/06aYFPikWC5pTmbk7QFcnAgaP9Q4/oOVM
QutTKq7YxYrFWaZH4IJ2neeVfvUs6bbFTKJEXW6BpsoL4mMD0e4g1P865ISv/4zS
DB9HlK7iGrIJRXL01XnMZpBSLC60iljwT3Aqk+W1RImleB2/URgUjxcw8SXTosFu
0Pa1KqAQouCRUe6nNC3uuwYbvAjTXDmIz/MIBVNG7qQ=
`protect END_PROTECTED
