`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y07TXFc2lzbdVtFHM3CmzmqO1awfo9V+3SxtuWgyRzHSzJed10RUOCdcdRQysSEM
K5YuuCbbnFwERZzUA3a3eo92XOFdrM9xVAOt0OHmmHA2K33UaCR6bsJLa+4uVukQ
RPRUTZYKE9N8FHTDn5eMu7oTCK9D6woVngh8j7aj136kinrEQt1wuGosly8+eoLV
dGkglICbVQ4vHFCYhQwKErtxjDY9oC205RIFxq8FxFhm95SbcENthhCmBaMDO7eW
c44Lo5ll9EWJA6WP7yBXylSOCwkX81+iq/u+59IrnCwCw28J0WMUOWfiMgzjQDzF
e6GrgGpa7rgSk3pbLk9EKvmhq+aF10vGO/dbMY/H0NLPNQnZZBxlN3TDL17KkZgS
D/DkNMpHi8GAH2cXjG01au/1adVYO9TGujmqtkxfPo5K5wof69Sj04HJ+duu9iWG
oZSle9tFAflKLsgyDaHzGI+DoXVtqZjQuB+gI/gjJDZIFY8xFRYifAN3JHz8nPd4
zQ21IRuHftcV8osVWMyfWASV0O3575SA6sV5daHqumySyYan+ieq+uY9YbajlJLf
7pjrj4fZf1up8ZmVVszirwsp1dh7ZRnDSnag3paBePgtSjtNlsIeGzWHyIxPKZnd
9Z1t20KXjQeZjhG96GjlmJ1q1YTGHaRTjLJqjD8rGiNEYIet2DWtN0EjwiBITjqA
hdYq2Pe8HF5fo2NjQMHXAwDg435ZhuulYjCvytPveXLF6bvFYzwmcgVAc0v8vPDr
E7na2wPZkyvZIwDA2VbP5seI+lkR1KlSdK99Ls06CNbL5ul5331Zlh8r7F8mbbGK
o8q7hhfQsqeK4RhZlmQbpcksPi15ghci7BZSly2YiLCFRPEwewSylMbnIIOPvQFh
43mAAg7TVE4EH4MVqigary8nyI3wy1Pr5JsrCfiE9EH5NJMwh53jcx76qItNL1/d
ejHz0jlS/l88vbQMGfQkwyslaH1VICO0HJJJTkLeioCWIJn1Nj94pxVTzPSmjwem
67t11x+qilxyoWEey78b0gVD85GNdDSG5M2KDdw67uLSydUoqfTRncFq5AgnfVdv
lNUADFtgmRgeokrRGmgmYcpWpaEbv1g43AgRptZSD/ALVkGaFbkinrF9HPO0hgOf
gbN/CZq9ZOMj5jteNRc07SDarPPGNJvY061TG4Eyj3fNWQhRgzQnZExVcSHUS1Pe
EVWb3ulJa7/C2S95eoy8P3ChgpGx9Vr3J+AtzYRjF/DcYMiu3sodRfnvMW9KZ8Wm
6cO4uIcncAJboHD5kvHc3k5DZbMT4xR6Xod3WwZM38fSn80cTbfdRWurjWYRKJ4e
bfo0XYGX0yq5fNI6grAKoRt+Haxorx0NKwEwnokvol/CPR3BeDbRVaYOrNtUyn8q
DE0Gn6mE0y8PznArBrhsqENrBB3GuNni/VFE66+VNWU8wOdVHAUYZSgQh3isDbx1
h5qFz+PBbRHYLcz3jNzWqsKZudrKH9p09i96et9WQQkRmm8i+NtDSpo0cN5oDxRV
e4/swcn332IQmpHhQGis2jBJ8PLDiPAyOBOYa5E9nK+9L9U+to0rVVj0C/sKfPsd
12Og99eQqq/EuRNQW9nPl0kdrksLK/dzZJZ9U+CwmZ7DrXm9gu9tj+7MawjHNzl+
pd/ZIIs27LNMLHmUHsgR7dotxTpuCgocofU88sqCO1xm7/zpKVxX3ZwlrCxCxzyB
j+4TLnD34uJkagzQ38F+KusmMGlHuWzRL8Rfjv9Fqn1ai8Ooj37OpX1tMy9G4aKJ
UfA4y+8HzQLjL18G64TCHuKfU2aMMCm9MqClMpXRwuqzM45HhEMT+5IyLZoLSYpM
NPaKy4B9al4WaryUGFS8AP9UeEsrN0JJZdEnquLg26ZhEPziPGwVrJCVkSIHJ/8p
gjdp58i44EhTMqU6vlgAgmS0jvY3XHmHlpOUG2VramJVimmDvqiyd5UV/1+ORppz
Jr9rokOsotORPIg340Dow0RDnsd09vAUerauGtqVMxnrpBWmKNQd7Xkq8aEMVlzQ
JwGosLPRoBJ78RGVlCbbJAr+fdzfGSjmSjdwIFLlhxFDm05gK5zgcYi+5GdRy9Dx
bn6viUc8M3PAMVZckj7zJEY7FYVgBMd0IAwm0/o8A93AVgooBs9kxYIxxaBmrKur
JMYFuHqlLOOBLB+ujyLNPym0tn16g6Xx7Bfpj0Wr8wEdHNHTZ2vHYfXSo+GWH9J1
dvc2ZZCB1NV3OptCeCvou7iixGjewfrmXO+lx2xZsuw4vpVJq925ul0HPPiohPCX
9ynzLr+g0C3uOkYi978fNWv6OdeUaG7oXR48mfr77BUw8ff1yCIlwACCu+Nh17cD
RlA5GovvJri2cbDoulY0hACXiUtnE1E08bqp/sV+s8y6qSo+rIWAJtMHzG07zfmk
RyDbgahf8HpNhrgjrU6hG7UQJ6zEj4dfGgLFtRPYXelARHu2z8TiQrGbGayLV2wt
wALM46Li4Xg/Jp1UmUniTDT+6cxSstAk5WhPf4lN38zPVMBet2P1K6fqgreWjqAf
z1P/bbIXOlGnHFFR9oL/eSOU2BiF/H6fDe/RYW6Flq2H6cOmYzqfQGwcGvEV1xOc
Afw6T4JSS5Roeh3yIiValgmjfhV2PptMFYSiJzIN/IsTypP4qUQa+r6gMKW/Aq5/
bYI4KX7lXhH+3rB+RyF6xJg+m986UMDy1IJQ5P4Y/SksC3atFIiZa/AsfGNa3Y81
xpUefPjCQa5MIUpWTL/jrBNdjE64SR2smlM50ohU2X8ju1vo/m538TrHvvBTfIqV
nX+yDQGy6Akvtfq8cas5XX2OtqtycRjWtF6qDuqfwMC3VcpN8nEFs4oQZGfOS40m
PZ2jaPS3PlugQojEcJq3rVp6bXxvFi7PqBe215+ah495BNw8Kh8u0nbDfc2KpvFc
HQE88fJXRBCgTDiS5VrzQ4O2atCr+uUiZShPP4o8ozLWBaPCm2JkQFoXCAr/pseU
m1lveB/V1ROYi4mwpa2RiYYul+1GPTw2eXAQqpcuecakT2mcX/2m8lVYu94Htrf7
PLQ6mhCjUTOAiRoyQ1KLpkM2kF8aCzyDuk3K+DKplEg8hafdudtC5Vfjqo9P60LP
RCyv3fhb1yeRqU53CJncX0OttNTHZRJ+VgXFNnoeLOeXNvQiuBzVfS8k7uNKfAwY
wDIhcKHbs/vB3MV09jgoYneqOpJQthGHkufQAMpMQQ/Kj8T1qN4YFq469zp1Ezmb
42pCgDzTmP3ggfG39rLupT7DNf7B2GQQslUjhF3yGFMMGuPcWTS6K6MK3ohtesVo
`protect END_PROTECTED
