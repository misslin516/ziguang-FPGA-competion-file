`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNaRzg/Y7WlXKB3Frqo2YKtDVXvOCpZZ0YagFlGt8PrMDTqUFdr9s24UvaK8SB+A
kkZZ3/1Cpsby3tWUdDyXQg1NuwWSJFO55O8rsY9Q3DKD2OnuXVGxNTtC7Pe1Fx14
yWwfWp5OUDCdJ7wnOtxSOCYl8XV2K85Tk/h6iReJQT2BWalJH+Cyg9GEOgzEY/az
n6Mlm3RsGx4WDJdzpJ+YIovq9+7BLbieNj6zSitnpQQmgDk/DsfsvlJwZVyIZqIn
iRsgigIrjJfNEqrXo2R9NQ8K65mrpWizvaOASzdwp8vxHJKdBrKblGERTaxh9SHz
G9H7NpVbVk4BIJtSVWTvfHfzOmoQSn9Qjr6aYDLy5rWIqLQffgKkTLdqXvB6yzWo
pW8asWXzv+Xs3M5NqlUXF1v2dj4qZffvk9ObvEAiIWwpXurqlPLilbBI5SB1EhRY
5epC/KlLiFWzMjthCkxasurAynyU/BOQAHIuyLFKc01hYjTqZgvGM2Lw4rAPLlYn
SSzU1+cR6QRL2bbNMqJSAbO8tPTRrjZnr9TjrCTpVbSu4Poj3K0yWovm3+b9zd6o
KmyR+QVMUklu6hRDDphiXQ17G5rvhPFrpVtxgJKqjtGuJdo8atVTDTqeG3Hur9/D
4GAZb/WU7TPrA8fu/g3bDOmtPWKHzqg4rZcI6hcmU1qwZ/xANnD3csGfOp9pePG2
EiTNGOz9zFj2bYbriLM34I8GAzXpgZhPpsczkLSKaF7ayr6wC7/nnA7IVUmQRa+m
6WlD3WDpbQwmN/waHcfOsw==
`protect END_PROTECTED
