`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/3rEEfltAMHckryEM6hq2oIhJ7+1i1lCy831LN2OxHmbAtgvORdSwYXcxeIJ9qz
y4a6HoW6g2HbgFdWtq4DXfJoVORBi2mnuDL1Cxp35wRlYhyaUwTscGr7+umo5/lo
pJTQvyOMgrPnTOvyv1JCu5v0aBjEwi0aAyH1Bomowni7lserE5wlk4RFChXJHefj
oqfsL4wV1Dqlyur9kF7m5cT/7IUoTUEQTfFEMreSTxk20mJKxH812Ql3BG71jY7A
m8JnHAIAwggCTlqhxe5yt6ZfMOS0wUCPrSBpPo/bhga65t2gAv7fUgifBGD1fyLL
67Um2SIBpl35oIzpXNVmzwgsqdWKK6u/QyuLOhHjHPm8KAp8SfPAdGh1kqxzajTR
YBBKoD8Y4bJmRCLN8I8u4eVGBejm/31ClavlwR7/RSqnTssn17LoeawPr3xbkCnv
RV3IgpS89xfwz3GgYvxKUUujMUE8u88/8tVDI0AUS3poCzrrjA7En9l+cly3veVE
Yhy4y8n/Kjxz/bcK2F1F2QetOq034Ox5tUk2euHTVP3IwBdece9GB8RiLBStpmTe
qSFzhtlVAIKd71RcXj+7ZCTPGQw57npW/QiWcU0toYE+TKO0tjzCfTv4L5eAUXvP
jRSZBbCuvUcCWFXG2YMrvqceXG/RZ3YcmLuK8VbANRMmTvi+qCpLdOcjBTPzsjKc
8mLmgIVEuaqnVyFh9ud1zB00+F6Rrl6gUXHlx6ABCYWNo3nLgDpgi27vb+ulX5qf
0jGtXPyGfWMhNBmUUpkwGeHOMowzgOFP6UyikvCyHgPERBbV14Kr7dWR4cVAQqM0
lf43rAT6xJRlT/g0QolMcrVxaJRxVvWjGmXTSilwxrQbTVbJjUV8D+Cmdup/uCLN
YwbOOPCfQBOuX0zmTZF7hTD6F2+4tBWCJKB/leZiMBDkWECtSnqw37cbnsbRg6Oi
6xeYy1OKQkjnymMHGVXuknWBVUVFCix6sWZqdqDY7EIpLTfdPq2ZCUOayFHbF6Wd
p86iKXkqDrKGGJTlRVs3IL32giLhwsrEUol0A3glk9w4/InGWS0446LTkhf0ag0W
LNINOfZvk3DOasPDLWiCfayga63jhyPI0V80wKf4afqvl8zdGyJNdMAyjc+rg8Xh
3B5eumj0PyPLwQ5rVdPE54LjV3CzxXfXV3hckxbzkp9aiGfDF70BJqFOVZAhmq7Y
df2PmnKmgxFk0NDwd+fRg07UOz7vj+qSweHtDsZWkqgJlevMcsX2ShHxmOzKUEnO
UqB1dXBt8/PlEoDygD1HaIUvzXPD/gdpTpcCzRSZZOEmuFhzzZ24esKu8+ctJcUZ
pwMWm4MqjxeK/CWuwYvpWDpnWp6ruTSJNBUXI9IvOmogGvujOlKmR9rlRJE/fjNO
q9iD7I170870I9EycdLQZv0fzu9DstFVnA11L/Pt9T+IJ7E//sFhklCrzkqxaUgA
SFYt1Cm8KNgMz8YuW5HTeeuB1Qe89CWbHHjw/2VxDqHELV88PKqHoH4YM6TzcBog
Uzqq/0MFMXYrdrQw1gNnB637qIFPzoJrLnVVXrA/A7FhpDerlcslhGlO7WurDvZo
qwKhEgEq/VsN40MyYxdpPGLwPCp/RdWieuop64pHgWvz11Hst6e3i9ed0yNfEM6t
p7p8ReNHFKtAisT3kE3S4l9YjbiK67E8ktnhuL513aTeeCh0EC6wTo8OTEH57y/+
33iRg4AMyKB/VRAuO0gY0JaRcxKymkKRsivPDss9g3Ul6ucF0iv/ApkjXH4thQMe
/++pmAtmRou6m6a2FTmQUg1yuAUn2WIOEzoUB7zNGwiTBGVWV4XKb0GfwkBpdnm4
70M8vPY/7esE1CtD5JmspHj4i0V2lXFwHv+FZbxXJfb5xQ9CNLZig3H94CfF9cg+
zMNYGQWBHtfJ73YoVfxleSXM5PlTCVr+mn8cHiPZEIAl0SflvZOyaZ81A9RrPZYY
PCfzptUMAwWzP07+/OZxKv7C/hatOpQ3CDfFWZYocPh8nIn72GP22YZWA87bwWVv
999m4GLHgtCT28vh0IW/oXAP2NVA7YWR0y8ONeHV52Jbo0lipYTBi1xplbMmDSzu
cDZ1//04eycRppcsKTdDwPZDUhkRvpQeKtKupPqA/2hCaZRFbE7q9+NebovgPZKo
0ZgHRxVAtRWT6AH8g71+8i1q6yBKDz1Hnl2ptT65++8Ftj8n4C7nYak691Acrz+E
lD+/d9TPj0LCCXOHg2+HsVDPOhSRA83CrRX9YYrW3XWqGhnS1Gpp7s9SI2u63ybM
8iZRuUt+lTosfIKdOwdy4e6bWKqRp/PhJ/tmx9aFzUHLrQeXlPk0B33eCtnGJ209
VQIO69iUXtoekj7buPQMv32O9mFThEl8/PPW1hVDPdkjZok+nhirZZcZJIhgj+9l
QKaLC+LYcxlnwfZu7QecsBELcNGOxi/kEkpXMG5iiwP8dtXahwNh9niYxH7yr+f6
SIRVaqqfaqnzkyQISelASws0MKxwbyCKSW5ZjcpNTmcKrxSMCg+dSTIloQddE4jB
UpP2vlvnd9BxaIVo13DPWkaxxvXuCuHIvkIVvTuYTeOvTNFiDhQYOmJ8HLYYOCyP
8OHI738Xp0kM8cZTISUMvKzqhVQQvVR8jM9hJToAY4bOWawnyCv5Zp/1aepRk9gQ
r4rpFLGdDiZ9STpbtp5KtVz3zFiyF89jwkP7AiTUTXmVz+/Zyq8XvNEFwzTg9MWQ
BLJrM3J/lpCms/CxN6Qxunx6EWCnGjZnl6iuFaVCrD2CPnCGHvcd/AatHTUnZfZ4
/O0cN3LFfb+J7jMPBJ+9HAafX8a7g5NFCNStCX1URhntQ3U/Fao65Yt5q+rIjl89
sJIDUMkBr/Nu2SNiBTPSUsfm2xxYQ+6bb0P7njTOlPQF0QI61B05kUNWYTneURmb
ljYCpctxUT5tcrlVOwyzTUl7Ib/+2xpCD4WJfVOGl2A4a0C/+Dwn5fmTKBLBnocH
XXKlTzxZFu8roy1Uyv85eDVJbbpMEnSeR6NrBhtFwrqY+pqiLhe5eLKDh2tDfJAR
tcc0S5juD26dri9S4qafZvNRfp/lp3xeDnSV3HYxJQLW8Fq6Aizg7ik5N+tEmnd5
C4mdHRoCLFsbP0xiX3EArbfv4YzmP8tlzDXYmbBRPUBeAPo+Wk1Yrz7Gy41OI2qn
ovDtTNfdkefytfhPGUBOKY/GAzRDBf0t1p3X/cmrhLjbugHiSdqNr6NFwugIySzx
7hbYNqLv8iwQxBfCya1jxTLePWpLVC3MpkFBtBSXB+FRk1iU2pQVmvlXRnegcyx5
iJYvJrgWDI7qrOiuRtOf4FIZdPdywzsnf60XsU/a6eiPY+zPd6eDd8VUc/H3cs5h
2IKpRJlowjRMbEs493x0AKvvgo/OmjvPTYFtxiiM/pjAxJj84ActCHZxn6tlSGGm
7Vpf3xsRZfJxbgUi4DIC8feBxJ1aN5Wn3SH5nVjXFDPujlLadMY4e6tIo3G4uuE1
jkgVXMoavjuh7EdmkNpvSJVhJuyDbOj5J7IXCLEOj6EQRKIxRhjw3DgjDEjyAJoP
Jl2KH00lgVTs8p0c5dIvKy4u9jBzY01YbxDcGq/U1+GzD8R/6S5YllHO8nFzYf0j
6GtAxHX6PKWMXt3uveaIcHZyUo0zkwxNQBPRkIzXOqdxBuBrq6OxbclEPtI7Gc+w
9we+9QJJBz2U3nc6yB5vBeojr889Zpnl7aEHSTwp3QNAKPvxjZJK7fMcSNTmR6eT
Ja7KaE4wZHvCunRYUMdEn6fgOnACh6d5mBRCXvoqXdZ5pKzu7IaMEuF3Q2f96k3v
tZEomCKg9nbHdPZLkZRTKRFP7Hg8EhN2nMJ0InM9KJf/krc2tBX4eZinQsFZOMgP
BXurSy013fxKb0BLh4zog6PHPhXCB/hQjpd/bgjylYgREl7b9FCq/FwF9eSi1bpz
HVr2D/nW7wMuIfgUHl8YNE6cJJBg/weZIm+FVLCcjbNxP1EHl5cFne45uMa1/hn6
Nf0IBi6sRaDmg57LhMneANj9Js1zOrDFvrXUJ9Islg5j5/fuXCyfctYa9LpBvMBF
b9k+J0T1DKkiIralE6VfhC1+k63MQh2jcV7k3aI9ZaERTo1yUUvx62yDvKAvYtXj
oLDpeZVLMkbdsFfi16uiEktGJTnqPQ2h5HTrNx0fgk4TNG+tkkHInpILjHNyXo+Y
bZkC2bZ6p/hOmO+4nIDKv7c53r+E7EAU6cwjhljfMrdrnut2Hz5aMEVrBMC9ex9n
hx46S388NbEDyc3rWTYBr1NWYTuJSc7DK54SanVLKu+GQjdXG/wT6eFIp3r2S6z8
xdUqnM+eHYOMmnsTWDTuCd4NHH8x+jBNcwjMQSTWN7jgFcdHC16W0aGX+0oGhGma
BxbmrIZXolQ8UvdIOgjxOKg2L9BrPcl5BUunDHAHnLqrxsKgwsn2GaKtEGpo5A3/
mFfFKf7W0W71CWsP2lZC+PjMYpYxoCByGw1HLRbVR0B7no0oceZc4G8xoBAbd4lL
m/iP3ybMT7bkZ3GhIzUSzhTBNdqEHD+w8N/vph6Lf1RhmXUbXCZqCN1cZAMO6DgD
OtJiXHOI2J1dOXivWFSCSacvG699OAq89W7dzqJNyA6GtnO9NCsTrm7Vwvxjpk3d
WEAFxRsjlMrMCnmFFCA6JE0edOu07hfhritA8dQxIYt08HbICtO7vLIXmjwoNhxU
6ScgdOjM5W8fFbaCbpU1iBJxGCvBjhoo/7p0CK6v98e7PHhgijZ+D9oJy/bObPfB
b3AORu264yLp3i7qDn3CbjL7OwTO6fSqSDfg1HRu3LsYts1Lq655pjOwEmMOyZ8w
`protect END_PROTECTED
