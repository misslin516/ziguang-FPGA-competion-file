`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mqCrDN40vpgzXz0lk7uUJXoBjZKpmy7q2S8Fl3DBjJ8+apJax+6FrSxfL722RDx
du9EKxDJAOZi99LP8B4u+1fGXn6E4LZDgNhO38Ic0H71bIPeyfYVw1EnN3rhmLMb
HIVtYV/lgKFv1tgiKz0/u2+r3jH8/xxFQp+4M2JbZYCCdezEoKcDguQhklj2cKrX
2FUWQJS0+quRlcRF/5kbb7mw8pdpBr7+UqGAHMF48LqSY69/0z3T2WjFFfQ6XN1p
pWYOJMhhPtSenfSkStTEuHgrHFIxjF8A3lsn5ab7F24bNmsVexvdrnLV+xKQ8Pxj
pOAsJVwKRPpN8YQdGedf7OfSupsFN0mLCSs1F0NKpV4C7yPFRlxJhkKsyozY2YUi
vPqLf/HtY++i0WirQj6WD3DqdfJ7TCmMQdXlTfOANAVLAmOlOc+3Kw1e8mAVn6X0
qOPnO+Dugp7Mw5Xe8kLwR4cc6L+1SkrZU+XUxpZ6eeJNz8x15MJNaDI+9pMwBlMN
pYn0nF1akoxuh+RjJGIhqbrTdHfql2KwG0GtxnfHAa3IDK3oH2mcZsuIQJqzlO/G
kzNyrN2ls8MO7F34xK4FgUjHywxOQ2cV5TX4tL95W+HRVHIpJ0ecQaSdORfbUnMt
zeQsUa24RRxHYkrBboRCGaqu5IgbAyLBFN/w4h2Bk6M4v2K/+yA8aBmF6Tl/DZtx
nsjQj2JtfaR0jyDuFQj6a7OWckE102Q26TdujnXR+Ay3BCKlZL1dzbxWr7HkzHbL
HfNG7jiSsrkH+eWfO1f0xg==
`protect END_PROTECTED
