library verilog;
use verilog.vl_types.all;
entity ipsxb_ddrphy_slice_top_v1_4 is
    generic(
        MEM_ADDR_WIDTH  : integer := 15;
        MEM_BANKADDR_WIDTH: integer := 3;
        MEM_DQ_WIDTH    : integer := 16;
        MEM_DQS_WIDTH   : integer := 2;
        MEM_DM_WIDTH    : integer := 2;
        DM_GROUP_EN     : integer := 0;
        WL_EXTEND       : string  := "FALSE"
    );
    port(
        mc_rl           : in     vl_logic_vector(4 downto 0);
        init_read_clk_ctrl: in     vl_logic_vector(1 downto 0);
        init_slip_step  : in     vl_logic_vector(3 downto 0);
        init_samp_position: in     vl_logic_vector(7 downto 0);
        ddrphy_clkin    : in     vl_logic;
        ddrphy_rst_n    : in     vl_logic;
        ddrphy_ioclk    : in     vl_logic_vector(8 downto 0);
        ddrphy_dqs_rst  : in     vl_logic;
        ddrphy_dqs_training_rstn: in     vl_logic;
        ddrphy_iodly_ctrl: in     vl_logic_vector(2 downto 0);
        ddrphy_wl_ctrl  : in     vl_logic_vector(2 downto 0);
        dqs_drift       : out    vl_logic_vector;
        wrlvl_dqs_req   : in     vl_logic;
        wrlvl_dqs_resp  : out    vl_logic;
        wrlvl_error     : out    vl_logic;
        man_wrlvl_dqs   : in     vl_logic;
        wrlvl_ck_dly_start_rst: out    vl_logic;
        logic_rstn      : in     vl_logic;
        force_ck_dly_en : in     vl_logic;
        force_ck_dly_set_bin: in     vl_logic_vector(7 downto 0);
        force_read_clk_ctrl: in     vl_logic;
        gatecal_start   : in     vl_logic;
        gate_check_pass : out    vl_logic;
        gate_adj_done   : out    vl_logic;
        gate_cal_error  : out    vl_logic;
        gate_move_en    : in     vl_logic;
        dqs_gate_update1: in     vl_logic;
        dqs_gate_update2: in     vl_logic;
        gate_update1_done: out    vl_logic;
        gate_update2_done: out    vl_logic;
        dqs_gate_check_falling: out    vl_logic;
        rddata_cal      : in     vl_logic;
        rddata_check_pass: out    vl_logic;
        read_cmd        : in     vl_logic_vector(3 downto 0);
        gate_check_error: out    vl_logic;
        force_samp_position: in     vl_logic;
        dll_step        : in     vl_logic_vector(7 downto 0);
        init_adj_rdel   : in     vl_logic;
        reinit_adj_rdel : in     vl_logic;
        adj_rdel_done   : out    vl_logic;
        rdel_calibration: in     vl_logic;
        rdel_calib_done : out    vl_logic;
        rdel_calib_error: out    vl_logic;
        rdel_move_en    : in     vl_logic;
        rdel_move_done  : out    vl_logic;
        read_valid      : out    vl_logic;
        o_read_data     : out    vl_logic_vector;
        ddrphy_read_valid: out    vl_logic_vector;
        phy_wrdata_en   : in     vl_logic_vector(3 downto 0);
        phy_wrdata_mask : in     vl_logic_vector;
        phy_wrdata      : in     vl_logic_vector;
        phy_cke         : in     vl_logic_vector(3 downto 0);
        phy_cs_n        : in     vl_logic_vector(3 downto 0);
        phy_ras_n       : in     vl_logic_vector(3 downto 0);
        phy_cas_n       : in     vl_logic_vector(3 downto 0);
        phy_we_n        : in     vl_logic_vector(3 downto 0);
        phy_addr        : in     vl_logic_vector;
        phy_ba          : in     vl_logic_vector;
        phy_odt         : in     vl_logic_vector(3 downto 0);
        phy_ck          : in     vl_logic_vector(3 downto 0);
        phy_rst         : in     vl_logic;
        mem_cs_n        : out    vl_logic;
        mem_rst_n       : out    vl_logic;
        mem_ck          : out    vl_logic;
        mem_ck_n        : out    vl_logic;
        mem_cke         : out    vl_logic;
        mem_ras_n       : out    vl_logic;
        mem_cas_n       : out    vl_logic;
        mem_we_n        : out    vl_logic;
        mem_odt         : out    vl_logic;
        mem_a           : out    vl_logic_vector;
        mem_ba          : out    vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        mem_dq          : inout  vl_logic_vector;
        mem_dm          : out    vl_logic_vector;
        debug_data      : out    vl_logic_vector;
        debug_slice_state: out    vl_logic_vector;
        ck_dly_set_bin  : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of MEM_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DM_GROUP_EN : constant is 1;
    attribute mti_svvh_generic_type of WL_EXTEND : constant is 1;
end ipsxb_ddrphy_slice_top_v1_4;
