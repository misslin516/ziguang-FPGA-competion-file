`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWZ6Y4ucazBRJTWmRbENHoaUKkqUBr/agns3yg2Xkb2pbJRBpyBdf749DTvnN0Wb
w2ZX5FXDKltaqXaEO7qPSo5i1zyJ3qYq25Q6EmEuTFgKHonrMi+kf9EmhGFD807X
d14wQUPapNS8WJXNGnC/DUOKCtu0r9kWOLgO+GY2mpAB9jF3QHGJh1v46v+EEnnu
OQ2F330KoPl1rHxIi7Bqwmu2e/ugccsQydY5B38FoL6ZeerG9LCq3vmp4vdKNDim
L6zgg5gbsd1okgiZMUkY4jNImEucGZ3ahU41xPjZx+iFajiHYJ/q7zKpJcxjrcun
VLONy3ppGrWNfBQreTsz8I80hLt8itlLTz9NxScrPAtwalF02X/YcveEBvsV3pgo
61By4jmrJJS4KKVSmZtpzG8Sig/aedN3NO0Uv6AUwGb4CWNm6qZ9StlIIBBKhF05
Y/0UKaODBuBGjXWchN5o0JVsUw7tTf9PCW8H+7QpZG3ZmGgOUashSUH1ucBZKnPO
fcTRdyar7k3GAui5c1MEV7bRcftXJD54W8OiFCY1klZ5VmR1ek/FxiL0cRr3mrI9
61qCBKpaLPvHM9N67rjQ9ICH1eHLhESnASRrnju0renCyC9wKxq3RROyVV5YQY6d
SDIRsEz/089EQl2dkVvwrQEYvVwYNh0pEheAWsPvbbnAijgSwfNLTpMJ2C4McVQk
lfBCjfCOExRDWn4RU98C5+5ugMspTe46mp5pdKMoZsmC8wB3MZ5shS066CaRCzqg
Ii7bD4H8SN7Wd8rhHuDIPUr7oIGZMv/DFI6Sx7ljYjcAkTsI92NFSo3YDa0bhV2y
nngRnoVU/LUcTJBYMRyP+SMOiBCiy36up1w+TWXSndNE+dvVVw1+bzV4/pR/8eHd
h1JZYUj6kDLMFznZObzPwofzNm1N9wxrYBrWW7RZKs3NJO+k5s6Bxrv77z/Kx4Px
6utjrt1kMJXz8zMzdG3Sg00IEiRWrpjKJP2JlFPv+Zt0APIb/yhsiChoJCHnJYvJ
Gip4pOiWxVWOq+lGsTNb/DlUMM3PQ/lBJOshHhDdAL+kUcYggFP+RjjXb+ip7t4c
yEnSVFz3u8+SBsB3kygGcPEjAQYOZPXCTp6GzzQAka4CZvsKaisJiqDK5J9pYgua
2RF5mymZlhgelPyC8O2uhXPXx+dxHw7MrTyM6Cda20Ck/I8Rkc98b6RLjrsBzCKq
lgl2mCSK2Gqxwwv2r3cDn+4WYKssYjPTf5j79s6k+WshWSwH0yyjKzN2HZDEGzOC
qUBZ6P9OT1OBwP/kzucrk8o6T4az81iixdIXvP0XJy+NfhSQNUotpsbhHUBQ+TPQ
VYV4a2X7F/BvPvyIC9Mx/6aXFRb9OF81Y1w5oGmplwVmlrQ4EDKAeMqOwKwxZ+wK
QOsfhEVVQFworz06CkOlBMHNlRM2sTl8Cueif0k08r+pDnyvg8uhXuis68TdU5GC
SaA0sE2UJZKSG/xifBGaBialMYpw+eqbHTCMogngr5SX6S6j+1PN6bWU8olr2QUy
K+O2C7BC4IUH4ttVL9ClkMqgBaYhVidD5WA6ajgs/pFQvZ/MYLsOU2R1bQkrGmwW
gRh8LSIBoXuIuWAkWpPYp+IaZjJjxiddjJMWLs6TMbw3E6J8LEcXrPiVy3NW4s5+
C/nBOWORlPZYwcYOJcWwqk36w55KKFw/r6wwPLsVbWDU7HKnjsRYEODLHXYzs7Y0
QzxAC38llMldQca+baWukeEMA4G5ocYQYmLWashRkEDKfppnJfNgCW0JEzjeN1X0
SqCkwz6ZN2u3L04DIM3PwOkEa4O0g4gKelYGF7hhbwQVBgP0LHfFJ/TRMMI4FGs0
/V+YUIG9tFFYGm6vaE9rTRTC4aVH9xezyDKIG5d+wjbJL/jPpfunAyw1fhjLbWyj
1wVy8gyBwrD+sI4LjIoP5SG3XxOGC/rzy+FuRitSsrT1rf1lBcT8/zy4gWRpxHiC
yUtw+iVEAjr2Ox8n3ps5uCy9i9IaKLhBY5FCZyu/N0SUrxXq2OajAIIkYZm20Fn5
9SVN0A7uz1lDIb+vXJ5acyyVRmQ1qXMfoVhkogrFH2iwUxyR8a3bdLrHQUIvm7+J
VFzQ3UHZ1jWpD4rWo8RH8wM3OQ/1c+Vy6qZ0ePHZ4rnV+YyemLqOp6rSE4ylD++4
TusmAnMEgdLgZ0btdSpsuw0SeI4nUYhyEaZHw/2hnVaCnpApb/AVcnJqNg7hdBXA
ouIkDZzox+Xii8BMI2dKkoMsvggfUXJb4hINDAGxv54z6APLi22Ni8vsApG+kAgb
`protect END_PROTECTED
