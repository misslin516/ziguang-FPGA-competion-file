`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/4S/StY6OOhFUcjsL9Af5Yb6WIiFIiRqUWXzYJeXECsPQgWlRQGWw2NJJ47Efop
cRu6075cas++e/dyxpBPgQwkMZPn/Gx28UsBdHUqlzfPua5yIIMIyjd09/Ur/fRT
1f4vPWRAq+WE6Uo3BpFA5p7McIUBvg0zxdvEWyGq+SmAAIN3K5HRhBmEcFv52oYF
ylDw2ns2dzKRaUY2gmCRNL2sWU0GKHCSFcLe9uiYALPu5AsDodRai+iIg8QGfNm8
hzJfZ2xC4QwOwtupmR4ow1eNmy++UoZsVkj/S1sae2/xiDAYpU32TiOi+7U6g7g4
fwXicZTWHU/YF4p6nTlNsIsyH45d8w0cmz3WZzRSm36WFZqx61BD+Bp4ARcCD4Qc
u3TzthWKZK7Hkr9YHdjvU9UWve624sULKRGufqwQBFuu7WGu+1KOkunPbWDz/Opv
5Yz6S3SFs0euETitZjd642vVuhdaYw7yncrz58H8+aUDXjB+Ji0/SfA6x5RnDJo9
DFB4FVMH1Lbw7OKb1PpfgAn7x6JYbLs3efzi/5rs8YdbGmfFbc8CkiY16oEPV5BF
xW8lCPnmphgEwcgnsnWDL1M5lXi+3HYVgDAM8tlkaoGIdb1WBjYfzOCugc9LJGJq
jN1imOIiPdcqhnNRHUX1xVkxWd6FCTJpRTMeAONsLIa7zxf29TEXLNwS4QDzAtqu
tkUsUfYlP9B4uk2JJ60674vpiG6N5+Z6LAiLp1r6AJwagiJF3CelGxqnsnSyKSqS
gAIwyn/QrL13J3nBscep7C+8lrxy0NlFARI3hUJFNJ3cY1cQwRpljA0LunUO+W8L
yvRWy/d1jeY8Nx088iIVYxBdKtkXAe0Qc3lCRoOF3P2ypukeTV6xo1Df6adIZq+L
3H4JRotuJ4Bi6CQ0gqvcUKzm62CKDX9OvmmynhgK65yN5JHea/VvqMupErtBoajG
`protect END_PROTECTED
