`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+NnHsKWRa3a4ahSxJ4LIdoLQ6U5KDBijfFGsYkc+bjtvcgPG5dM3EQBmjFcy588U
PUcWKCrrdbUh65u+sUG4cqjfQMAHO+H54cteKadIjJExHzxHx9IzkFCtg3UmoMh/
bWhbpayq+erzsnljEvPBPsnwoVGcIJUyEDgKC3EMTqo1fAUl3LXpsg0SCOVIVx0q
FKhe/wUHYIzYjywn0PayduRrTh4D/qAp6N+HHxOp8gBmY46BRY/ebaIIJbChNxpA
aTRaDO62BQHJU75HS4BWGKUwNb7gOcic8AokK0RbrPnoDOy2zuLD5X0yMmQU9jJ4
kUqELCFg8LQ1FLAC9EV+XdAI0CakSYdz0NZoLus5072CyHh8Lf1DW3E0YwlcHwX8
kXZm0YEOCRRIGnoS0L5dMd6KCQ8emRjC9jFpFx56P+M6mrhr1jGviioWZV/oQFZU
X+O087F9uSCohl1tB4lzxzVsg951tekYyLQHKYQbW+sINZ03A8DzaXNwDKT0F2E2
foTBHgUkh2eH70bCF5a4IQhqX3IDLaEIAdQiJ3of/lFN9L/tot/sJN5XO+tSOCtv
fFHcZG5o2h+zF+3qTyu9fM3Kt/LwkuVLc5No6GZmUdoO+lhDOGvO3Mj4Ly1o6nUn
M3nrDoO3Y8b42GXGZnwnttsEZGBUXun/io+K+5HyLuDE0u3QORXvC302JyEP+IxQ
qo9mnb+p64oD+HpbMIG2LwT43PSPhYMQtFhHue3RJsppmFh5p9wsEiZmHL2fTKMn
ZLSmt0/zmiWsfEXnloBOTr6SuS4sKz7HDwm9k88Q6Snk/zlFt+f0orqkOVwr4XWt
iM8ENNCH2ISTGi9zB/qR4++5uBuWC591L0bYjsBykDOsxzGNsiUbTyTPi0fjySdf
9LausJ5QgFbeNYVpF26MMhyJnUlP18wd5M9w4hj8l8dhewL3Dv3ivsMxlR5JhHcx
jNeFoiJS6ptR0SUXmbE6zCG6WKHK9mCxDiu8mS5usIDQEnqf7pnVSpE8YTYHtel8
BSztJr+QfBF/M8hapaZ7GTL2XCv2jy+yYPy6lV9D2iJA0zmM4sbLY9fVH/8inq7P
nLr7x95F0Im0YnITbLWtz3SnVNbS1QpocOWgor7GEhxEToBKWM5BzFZQOigV6n1t
67l4nE3KrE3qxtduSdKxa3auJ2mpbKzgKd1J2bcdFLx0dAia9NfIi0IIrFZViI/E
6141GQXOjD2sJQADc6ToTtELTyKJdnSg5XIP8TdcRSVK9JXIcehtWOM/9cutSkQT
czdhUDb5s98okvghM4/criL3okpa9yMoza8havwtthdWpp0NgDoyU5p7kISSa5tD
4fjgpozrnG5i1Oo5eDasZ/bG6HmlIo2hZE6MTKdWAQpAUJADd8RaGpu89oZ7fzWr
Q4NbGHSa8DDFBVSwbm8gjxvfRsjAfhgb6MpR3kajGXVe3W3Hs4gP27VufI5RqZo2
/3iMLi76fUXd66saXZ75KlhHpl8Aft8iV5hpX8m0lUiOHiQ7e0saIh/d/GoCdHHe
zftQ7/mVRBDjHsaNzzhVrYjDt0/os+wGgvvkdfXqJ1kbyXWh49qz1CpLZlveUken
3a8k23eNi2do51mf4OVl02jYu0KmbaUt8i3V+BgI4BXkiCfePWh1rZAPCI4P8t7B
YX7cnUf8JcQlxkheq79+Z//bihhRPeAonXSSIpXg0uldIuxUUnAadb5alhmpD5+o
ykoHZDoPB6vpWceMi4saYf8H3HMd0APoxV51md0VAHKCz+rFpvkU43yDxpTO+AcA
qgUFnuzj0LAvvYVt96ZlTa1AaRh3EwlPZN4qoPjQrgMmyubY/GaVzxE1P3s3rGCL
E2rTO2BMWcOGsThj9+DY4fcRFEI1krNAw/ht5r1YANBoMgZoqGA7ciFYINU5dYTQ
KolzR9G1MHF9f83So81J3SHIl5ve5cWwb4fTNFGUqSTFuv/hN/yTrSYWc6KVnmxZ
WEttLr8T7z7l//XPbGBRPZVsYu7zdVtrA11Uq8EE5auzOcBIo7iUQT35HtmRGVLB
PTQ618gmxPKjijAt9uMiEF0vSp8lIiihwz8vJbsjbNi10gw20buTtfpTeI/U16MU
YpqyeuUtJ2t0K4tc8sjtAeKeIH0OJcRPE+180yCsk7YsAFjfNvBAdw2EnLib7c5C
UC6tpaR6kFrjI1UsYx6xuOvTY4STjb5tfHfIjLBC5tM5C6hwbj4huSZ3eZA/9APQ
bOGrVR65PbRSeiNGCrkAvvdCbBT0hmfTgyrCb44dim508d3l7LcX9l2aI3EeeUYx
1sNdYwyjLPvdYpfINBr5N5J3cVWOZiGiTfHakI3kloeifwoFYdfJS9xS6hDi2OrP
9ohV8M32cyRgUg8EbQVLODC1ZDaKHZNMw7KUJKgVtwQuCO4u2wAGN+phe5Qi/o/e
Id3de2AoDEWXFKwsNYSb6Y1CMhknHLyPCtdTPtVYGbEMTHKRNS3OqM5CwAaB8+78
ebnmUCppEUgr+OAW7p9k4uTmvrN0FfrHyo5BENt69ZtjrQK1pQSGyxJl7zqHnptn
Wgt8eYlRcDd+7jAjl8WoWOAFDgQ0gmQmtTcSLwJ/Ai1yehSNLH/NUGxSsu1w/odb
k0/CQrFJgWSfOb1aOhoQnz97oDf5u8YIzKzTSUlVT92Mut3eFdMDjbSqgXi61Vbe
BcSGuqDFOVFqCjcmEsqBJ53+dWAaENKlusUhJltdRi0M6PYVfkiVUyN1ovHN1LeI
9qzdetE4bE7kvMg0th4BzlH18Gp0nUotD50sAyZkLfnZ31cIQmDATzxK3caOy5j3
hH//LppcbYsoimnyWiFNNVb6RPFQlvyfVxJT/iVrAyaUzoa4UV5uWuMrNv2cQWIo
UOsRCaF3oc/AgOVKkvXtezSb2g5rmOHv9p8sniXstWUfXZSiTX2ZqnC36Yz4sFFm
pq2GJWwRptGnHeqVKhWyjd5Ly3kYAG+DMV4XGhPbT/R85FVpxPncut+Zb89jNAza
gXTrAkmc0/EUA/bTsdCkfEgcGKpKoM638JLtjt8hQ5r0UHHF5oUZjoYoIHnnNm9K
prXrtMKhz1yX8SxDuvU2SAzc2gqNqNamNNTQkacgjsSIF/go9cOSkkpl/6DVKzqy
5YL0LKVx2ZYOqk50LhSmBbGAAObCO6w5A2kF8ETxhyspkklMCQE8MsXYGKW4R/8c
Pvv3Me/Sta9UMKbX2XLxFM1aqDz3AZIY/A/9wQHeGc//mx1tQGD6h5dv5u0WpLRR
MkTt9CunW7WFNtmaVOFnFkbgAfYyIoOwmav3pGWfaMDA7chCq5HcFASrfR+2rsKz
ycsTSKp/Q6yeZoUNgcG8ihvdk4EQInkfke5c2FRYwkcxZbQJQ1HBlos+s7AWjatY
tVvIYMdxuZUpX/2v0CK3KjjRdeW+1exwJ8bCV1N1I6ur0RuOFg65IIuJk/PNs4gM
bZebxxKT/7nM4K8Dlq4UdVt37C/4S0JKnEsONraur5CX+nqvjvrkG2bn/BY2LXcU
YrEwoZpoENa35t38HnkGfSK+nWT9jZKXa6Rr3ufivTecV4VUhXLx7/LhoN+zemC8
+KAka0yRz8qGbUNe3HAMl1cYeHXjkmD//foz29P5doSyLqrfjDMTuaJ/Ku10W9Cm
BTDE2+Suk4l6vEGx4RapwKcph8wri0pgbCOjFAF4r12yqG6kPG8GuGu6NHT6IVNz
KCX0NvVWfL+7iAq2qJOVPdirqHkbx8uIPwRDEpbLtdU1N4hdZahAeyNHbF1qGbLl
iXccwzjwmhLlE/QBXjWJSluELauS5POZeAeHu96N77AUzMsnvyE7AmbE/8hV9oK4
eirlu3J8fH84PFhowoDEew9xXSGQ6AmLp9G+gmrG8eJLQIysJf1yuSZfvxT06P8W
eVOm6YLVBAnLyLTeKcVEHfuJ7JZaFX3zwHV7ENEEJi9xPyUpB488J13OBdQsQuf8
206zIH0+ZZyBI/OQXa6uyVOdrWYeFaka3D9YSFOJtB+xVaBOkS+PHvkuiA5t38oG
89qPeNIgQv5r1GvXnhQVkyDbxKfXzAzs0/plWhivPiByjMobUVVYgTRf+FLo8MnY
asgm0ZPe0QXm9d8Oi+5jSIKjlFgFnlX/an9uG4JkCJQF6rUBSjVxtgqCr7nSUh5q
DmUT4Ef2UKuFe43/xG6yVMcOE/n1PnMoIT+4pb7hhhfAJvhJAGNgvUsi4wLZD5Bq
Lts1X//BbLgaAeBrmANukZlmYawEuvkau4BloST1BVyMuXWqexhzkEhxHlm5Oi9U
d42M5GPh6Cp3ThTJq2spbeMZ+I3br3aKeHKh7cLCmgo6mjrKyP2+fQm9n19y1sUT
VXmplRgecVzDDr4/3NZF69s7q0rIZJcuXX9IrPJzfQcS/wqYsSxC+dWBjmwT1Afo
6QPd94yE0AzXVYD1mItLHvi9nRhHVz1A2fi1eJzJj31NFdvm0qGhsLelScq4qSs4
M4qZPhDDpkf+vaHhTUzBA6EfujhnmZm2mqz+17JNJAs0i3qYYAWEBoaOSpjm3dxX
L0CgLEIOhLfyqFQQQLO6H/7LAYFCeAHgCb0Ya0Mg7xCsToQ3LZLqH/OsHYfrJkXV
GgmH+F/Xttb6W5SMWyCKup7MnIkFd67Fnj6DHtP5HiiFEblG8+IX6iMZT3DyZNi6
HFhb7X53pWdM5EXJHJu4r+AsPxbyVDzbZKavZWGpsF2Bm6TLZPu1bkxeDoj3iQ2l
Ys6ftA+JpM1DJ4+gvDP+hWlEoaCeO75arLcRXLnKF7I=
`protect END_PROTECTED
