`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kDi3Wcqn5LMK6leVih+dvmmS26InayYWvDVSaKbIFu/+Lkqe1p5AeQl7HVrWAx70
nW0MF6nv8pRqvySSIGGsPzkrbVfQHT+0PP2QdVojMJpiwdIVRS8gBaGKVTU8oc3g
k6x0ULmABnhA8QsWCJ0Z09j6LmPBaWPI8eeQYYcRthBuw/ZN4hMBITsupSR+50j5
Lxfq1ZDQ/hOeN2I2OIuJAo9te4KULErx3Xay8zoCNZn02BhdKzmXA8b457EBoTfV
xmiAZt6t7d2SdoaKHkLsomIuejhI6I+EEoRP74WTDzi35FNvi/PERQUUaG3kFqDz
R2I0BOLPVon5d89pM2MdUdwg+VcWHHTNlzntLYsH7YvhF+xmBzJBbigjbSc6DsxP
soz7jMY4fJhY7hhN1BYhn1Sz4V+NB2rOCyIcfNFbTdtCj50H6aEWYVALJAdeaBUQ
mPua3Q3v4CztwQ2EFnzuap4jTJlaKAuYfm3h3EKp8zuEpDy9PHzA/CqVPOIjQFLv
W2yeJirCOqsESe6hzsR8QULcObaH/+P++rsca/Za0wjvlm4zFFmfJxI/lQlXra1D
BMZzf4uZcVzkWRgdQkylPoY3/d5ogqlcYSuyYsmaaDJOm7DhvKWtWfvx4V7Cc/Vv
MqUxrUrkDuCgS1zRhKp4RILixDksA4pUhAJ3cl2LNmZa6UsaNnxhNU7X0rXM6l+N
0AiNNRa5634ErKDcwq0XZVqWUQ14mAynsL5gkMcl23Lnt0DB4DbhvrULZS99C4dB
FxfgtTfyZxGja9iQ5BMWz71JYYV6P1354/GnNwao5tAe1NMv32EJR7JnQVRAAbcE
Jc3DdGRVjkBYloGLgsRE5jcw0VUQ/2FSgE4gcWRQ/QCC1GAmXeRfqPsSdtG6vKRK
RgjnpbDolA7aIiFYuFid31+luALb+QvCRHy3PnDic11HYChC4TNUivlUhOrsG3IM
aJ5WG9dBuA0xyzoCU8I/Ttz/RNJXdqTYm61lcDcym4WZmT+NAgdHxuIfsd3nyV2e
uBBF/q5ilitH9rCs76uNuRwuDs9E4VO51uPFEp/q3r9w+20/0S+gFc4yXgCi+8Dy
LbxfsLrZpquqWdh48a7rYiMZNbqWJu+Z+vrKRvZh2z+9r+JLuSDTCqxggh9GDGtM
ro8WhVmH47nMMRYxypxn9WS1Pevk8G0HjDMYiyAFwCROPKCX7pGgvJ095cMXiyjy
UM6CXsxA8PlmIBKtvt2aIwGgYBOhINZkw/M17xmtXiyRFf08F9iA+cOHUtw+AMK5
nRCttf2tTrlxyNXrB5eDqdr6vWn5lYvdbBFywBd1BQw=
`protect END_PROTECTED
