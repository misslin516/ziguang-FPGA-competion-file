`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pa1KbFJoItLocT6dYFf0gqd7bw58JudAxsU+RColxYoErQIj17nY0RGtJPZvU2s/
1ZoJR8ZpdRfbj0WDkiCmPJs1ruxgP/DvVK+yKnSPpdMLpfGY0Ss3iufjaSX7iGCY
kCuW4kt1KR11YXkn/6E4GjWDR+KkF8KcCCzKhtqx/QaDI/bUkYfUDrkgkzBM7EMA
FOjMzRweOj4SGp+ROMr/FWH4Ri0U6ErZ2BZ6NUnUeCBDmqNMMFIZuElBT0HSfyji
/kU6RGDoUsu9vOr27GDJisNX4nIk8CrPR3IMCfuHh4F5MLh2fnV96DxRd5wwm00w
NzKBwW3nV3utW0lVS7SbOTifOuKoI5DTonqeEw0ebQNXZlpOfilDH/7i3SoT1TTn
yeH7Wx+vM/jaSaBeho/HpSB5H9t73xS896XGiPUlBOC1H9b/YQY6kozfHg/WG633
TNq1L3qLdoqYHArWP8+XtqO9UtJRKEvMhz2g3QBoD3lU44fnfvqdJXhw9htAlyQ2
njXcnBvbfj3RGh9JuZ+OKVHJX7BFGsUnNiXwc7wiaaWu1OhX2BZ6FlHVhzsdESjZ
fW1WwiP8ftnd9YltJzCCRAt/Qtc2Ki+quAXzix/ZkR3XrEMJik4Jxp3TC9IxfkrG
eU+slNPexRhuaFABLo7S9xzjOdfltlQ8eEvMnjfHOVF8XsvPSigkbdsfQegWARqZ
/VKlxuYokl2/4klSB/uPNPvotr9TkQC+FX8chbgxAhoaGqMTGGTZ5GOMX8qisJXC
mKW2SWwR9O0GVfRe6RXC3tNoVqOXdhd8gXMDxJXEKHiMH2IhsZjXPc4YZYC0smZU
OK1UigXLYb8rw2hbtsZvO+8TtK4INq3/DikLg+BuvpT+EWJ+sMO1y9Q8dw5Dkdkr
vQUGq5pJdhJMANZ2n3saOPAXHTSaMf0u+X1BE7q3pccWWtlBupJwP8bxoJUHEXgL
5k9tdVH69nZbUOgrzdfXFA2RJjG2YuWt7TaJ/dcZVTZXuhLgug2WXWBQUid4Om5Z
V+cR8dZs/TDhcxOdUa3aNUgLBSqESH19kXu8cbEB1Bwf7xxs9J9vsXf5ZyaViMXc
BCKVJi668PpfYKol0WsWhMTopTQECLht/cjrZMK9ZSp1vTSIjiMrNt4iHOpNWpaj
UOG905HFGKRJst+qwcMk4iiELsmiTUzPpNExYwfiEJnr4P62qBqTUP25vNtJC1fk
SpKLVOLD6e0RvJzk3w3F+A==
`protect END_PROTECTED
