`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ho73pfkWBoE5gOeNZbnsnB8b0vgIwVyqawLfSwfhR73qreKslqdqIa221ATpPtQ2
Z3DEnVFy7SdtrrOt6pZXdOX0oO4X6H05ai8TXz2OgJZpUllz1J20A8TtMCpBJY9v
sgRbFEmogFGq1ErHhIxTluVBB51BAPEN17FG8yBfRtv/OBtX24YYeB70rcK9xjIq
2l2KjIKhWHfNlZpTteZbtdyQB/fdoPG14dU+nBPx/ogmvLPFrUGTksAlN3u/VqJQ
ixDDGIXS3Dv9e+o08Z0uUCtWXgqim6HQKH/URS4dUEb8w9kEuK2L0Ibopwo/QESV
iFwg5JasS8oTQGv3WQ5PDfbmcaz9PNSnzjR2ueHgJY8tlbomxlfBzDtvBaASXXwQ
Z6InaCNJciLb25UiBnyuKbJ64K2Fqf1l2pzQEessgzY4gUT67hjBg/AITCqD1Dfp
5yRR7qrTsnG5kWK/y7HORBmYnXRyq3n5dIAZ3jZ/bKgvFmvNb8i/Fy6EJq8nN2b6
igyv0ZY3Juh97/pH+FyRXIz3PgXLKPv3cuQ0/aYcD9h6lZGx1OFPuCZtl8TGKrE4
IhovloNbnu0/YF7OkEVb0sIJEr4Fx3hywC+y3v18mKXdkNG865cborS5ue5UfUML
NghDnf/ai7DSqW7wsuW2Y0vOXFwQQM3xx3Gz9o30eCoXL308VCkh6QD2Th4B8eip
WVpU/chpTZNf5gHA1RNfbc8WHX2SS7EdbHGW2GQIrJIl1SGT/UCcAeK4uTBSvj82
7eQx7ZY5dlliGUUG9ScMMcL31Wtd+dsMaKJa0Q9U5J1Avk1EIAfed5LsfTNrW9oT
G3zzlTzDIRChpYpxWOhbbi5I4IG3/ubUDwyGfamdeWjVRbJ/RYtHQUZRYVmZxEkY
lD7n7TBKVXaM31uf2iPYkY8qdwjq0F5BI6vksEQQCkEu2fz/Op1X/RMqZh2x2Sqk
rGmMiRjAetXUhfbYhxKd/lBcOGfabGYUJTz4V95D8JeNlZiFe3E8rh7ph0wn6Um1
HHDnYFPVj47XBEfqHpAumAImASi+4eL1l3mnGuw/Vijvb2/3+Ec0YeCU9CwQnILh
0mHq3TVLXzwTPFa835lu7s7N2+eZKT2n9UbMbBTs002IcExTWXGlCz3BFfHrsAd2
IrQabuUu+yii+2cB9+YbR4tkx99Eir0xub4Kv3PiwrYjl4u1F/pxkyto74Jr8ZRG
3LISqZ40fwBZXmUWRuc2I2JaqdRe6e1i12RNRuJMo+shDNm6G9mP3a5kB4zOojig
6zQoDB8ZFbTqHJNeLsQnUzCWzyv4r+r/ftof5x9jRFKJD3qqCTN2Ynutjnm+Tzz6
ySu2Fl0bhof5iSlqmHkVgGFXDnyynyP6eBQSxWSFHrnXei3mHuJhvhfjyFxxOPWv
Z77BfXa7JGD3lmkzYpdF/P2JNbsxxjFqrK22icQK/yaYwlV9FBD7gNf0MU/wxNLc
Vdz84MAACrPD2LyDRevzbBBSPnI4mYLZD6I/cNj1boAYyG2qjflbEm4dVKoz8Bxl
2pxL8SMAoEcirWM2BELyprgQBrqrl9y6JeAFuSfU6wA=
`protect END_PROTECTED
