`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
778I4ICKN1sXPuaH3h+RoWJG1VZycMKZkhQvahyL37LS6WJvrO4PqyU/AjJPAE8c
MdTi2ixDujndAESG1qKx2AHhzehs3aAc2SIKg01osbhPvmEFw4okZcplw8RyI8og
UuwTrJnlStMwjwa68Vjxg1QzfMJeIEIOAVFYXh35wjBx5HfKUBbdxe/LH2NKJe4e
ZejUS+vrlqovNBfG7z+pw8MNoMy8KPukrE8/B67o1aeMRBKGx9bGbqZadwNv8obp
ahJ+Sff/MUyhbl00/RwHEcU8GUwNbpJCFZJoBZ6PHRpzZpG0B9iZzLypmCAnU5sU
EgH/1vad9Ji4Q3tGTBBnkudypVmhTwaQbl/+A6gOe6G9tnHEjAZ5QduGRAtXUR8m
OOgpZv/+WGtNyf7aGVtHgCxNDVj8AtbzTM4A4BG9Co3Ww/sZ/9OxWU8d917hGWpy
yo8rrJv60GuXVbz6plpHdbn/J3Uxw9YiI/XJX8Sg9uz1Y5wvHLp2an6vejRQhwLP
48ec1c+s7upxN56VJGpZKsuW/E9ue/22KaJkKVs/DIsk86Y9qxG5fsCfA499k6I5
mBH+5fz37TgcLQb21DV/H6zwE4aBkvvurP46FcSagmJDk/RziptRktD/UJ9xINy7
flpw6nej1kxz22q738kJkEaUX60KGR1yTI3f8Mfg1wlFXFZ5ZYGGccvJz9DHT0Pz
CCPA50t4N/GjB2x8rqV4hW3R/HUXDHM1YLw7ApQFZq51FKXBsEue9kq81SOgD60+
/wK6XWG6d1yKi1fUuu2tgIPVrXPi0+yuWApPDpHr2giks4ZPvQmIKOVJygV3et0O
XOED4oogxG5jKAYp5R2RjQrCt48YDmtSD1TgJCIZG80j+whG35e6DW1Ot1IGqKA6
I+dw4qaMvBfR8oK11ZIFbitXpahiIZ46ty3mfSrTKjTP7c6SFFJaRB5Jqy9nSXyw
W4SkQ2rdDyNaEN/NYVZv1stkZQZxT7y6JT/JewICPrJeyLxx187eUiRu0pojNn4W
qtJiHmQIyScQRyQ+EPrU0GjP4GUfKVzz8vn+Bqd7frmLqoEbBxhKXwx9fOJHiU+N
uokdXEAOCOHKeVgnBqU2Z4Pqj/CqgLwllGZI9PNHmZqolYAIZb14hRps1t+Nah0g
hSFdRm1NbP/7ItFIxC2FRXVb+Umg2mA1Ar076bxBzA2PYCr5L83RK6Gy7m0T2lp3
/2acXESUjm/k5ydDTtI1EL2936dWP/ytPxMOK/K7duzJi+eCv80Eo+qeFWH2rW25
QrF5npRivD/Db80xRRQigT2Zkjaycnoy7PAi5OtXhXRZqahpJ11yFnxrTIvLgGvt
ZQnHIFPHEaM+G82bNfjB+a9xHxwNJB6D7bIc47sVSbqOHwi7XbSf3wv/j6ji+zp3
kLeR3yzVsjcrmDi49l3Eh+f3jwwTHLZGhd6T15wug70SW2oJxYyhj8yTDuEQWcwT
xqmbE4rBt+ZFAN9ifjqdS4SUpL1CI0vAQi9ngAxgRYMSrJD1PF3wtTwX7yieqB0I
CYrtR38hf1shalyUclDAtdMIi1hKn99QAbCYx6kWZx/S10iwIxN6+FF1zYrkKCsI
W7CF5zv3R1ktcZTh4e+nKfjU6bsb0nZlbhSEFHeAMzhMlVmwVBUySqOZLikbF/LR
KDV2RB/PkqX5dSWIYPSoIRgtZmgkdnVEO1aeo/1Ak7f6ROE3HuDYbrSDjgq3cm5R
wXZYqlqFs2nlXYI5/aQcPAn7IfDc7oTbwTlceFtkVzGP+GUAidOnXUAmVhznZXxZ
+XQ6fG0UR4BhFLmHh9BSwO01Ut+g9dBi+/1B/jJFhOgOAFseEq5EAAbQBzLJAdJG
h4oKkSTWZ0RX+ZCFnV5IBk7iveKI/C7U05vbqKL+96baVaWtpc5YBR5OCdkx3Biq
xWWvtsl9hiA1BLItw7NjQDkERSV45zcuFTU2YMJBuqadIiqQe4W2NgnOOrPFMqlJ
yKFphLCXJHRxYWW/227PlB51HbeX7Kk7X3JvU+a67g+sOk4MsOIVxnOvxsdA2sYI
C1zRLANKdDpL1/SpDHTdQvjbJhvjhILkEfRpdfouRKHvN8Ee1qhQK7C/n7lGGDfE
0GT+ndChRPwbhszTlppaODIKhfndyxU5M3je/QFL5UcKHPYlbRx7jg+wCJ0Fyt2e
BH1eyLBUryj1IayzTBCPTLN9u+sqCj+gezMhQiCvBzW1s33NaxgrMKUtwH2iIxRl
FAtMEh54QF+Qm3wp4X8kV9s2NgjtFjwC6sR+OhhDUXS+8b9Ya3MR/uwsG7BpxLaC
0UNlVpoG2QkXXtbNHmB/4jsD0JmU81JZOcUPIb+O80752yzcs8KNOufhp47AO0Ao
qsd8pZHYkELrBS2iq0tLV0nHrsj+x+0WjGhnkeaxqB4/4kieutBYh5S9W6rT4kzL
W3mIrkybOjuTAiTrwK8I93w+7WbMG6X5u1b+DvRfQ+/qocsiU+9RDydo69jVhDPb
Zpw665EhIypPXgzQwFqV5Gb2QPFt+UahNa6jHViIO6nrJuRC7k5BEE1ZajV8BVe9
W6T1VMV6l2hleHjrJ+yaWqCWxHgXjwWdnUMPuomkUF44cT1/ZQrsWzGhozOgOemh
wfFhCFj+p5btQG0bqtdB6UanYMUqSPgU+g4DbNKTUW2O4ptouqvGXCAt/F5b6TZB
1bHyoL0rJ9Y8/btD/P9LbXLyTR92AGNowrJp1nAjwt6v6Y70tOyXxeIiggYmyZO/
IWrB7W6Y9GfVntu7HPETcILMXdbZQrmfGSxyFA5vn8aizu5d45DGm8NJX/olnGR0
TsxW/fglkpIgmU3KnmnN1LcO+7B0+vduJWhlzPdE2qXlVV4Glzry3hg1J3YP164R
DPJdRBEm3HbbMGXnF4hzS0qbYBUo3y8KiLN56LYxxMkUTzYgU4TULEsCF0GUyat6
hBhHChvBUwr592kwzz3fRYK+oLqcohJ2eUAe0lt4ohUnr++N5vOKbAlII8CIbnBj
4gtDsC9ENM158kRVVCOCWLm5zals4FW4ewX1D35PUh/W4rMUc3XWbEnwLHoiOYxi
s8BpGjsebtCNrCq2eqccJAFqBMw8vqzCDLmct9mkufyGT3LBxwvsHDOh1yRswOi/
SPjMvIGGcPvQwD8xWMnPYyuoVZktfTN7lAv0oBc17zQP80Gul9FTNZqkU1YdYVnY
AYn9K6ORpHIKSCRTN6Mu4WrNs/EEXfJUaVjebwDX0h+gYnXDF5+vNddX9fI10ONL
NK4QAKg0hzQYXNfA1vKzy2w9txjVjqF9eR9nhoC/siv2MhzVhWNs8WiNWfOeu3Ny
Ev2nuWmTBR/cd9RiUReaBtol25iRieLtxmY9gmsOXEsHGOuRTdA/vK9ayZrQTZN2
4uSWO234bLrEara0ZXRuq5UveIibCVrIKpSid8KBOWiKUS8ACXSvF+OCmyAvweHQ
vpyEghmhBAGLnrkZ2lwCijxB8RYFiyS7ab2y4UjManKj3Qj6TesJrYUdfUpN5cGj
KbZGbyp/06VmL7LSATxtTteOxMa35N7ao4HK1itkztpePtLvErNfqgxhDpNpMFtF
mpiIB+Iljiy20h4X3kc8dK1HjuzBa1MlqvWvf2mMKjEzojhE6pGrV8KuZdpA2Uh0
JZ5VgMpBee9zIzHP6+sWbvTi2LoB9KAfDSWFcxazHN4q5RtMS+26F1ulfqH65jSy
gecuxDb79FIDp5d9k/hKnfb4jZfGPCPscYBpS/z6Y1X6Z8JiGyUo+gIPqQJg7+Rk
Z04tJgJQ9y/ECCtgLVPs0u5vUjFc8fb0wH7c05qpZC66jJxwuHe11ziAVaEVMEUu
hF0BaecORZA6PYZ3SJ9pma3qh6ZAkCfZ0g6bRZX8BC5bp445O6XFHDQs/NbYbrjN
FOHEXI2XP/h8Ljmtwcx/CbO40QTKxP7kDIzG+Kujkv39tZEg5uxbdKRkKZ/dGgYh
QwwFi519R7hwwaI0LclVWlGm+Xwuo2HXkjpGpgN6u4pmdOUzj76aYfsNlOWiByNr
UNaFSUtoWA3j66G4KHBqJBxE//SsMsvS+J0ktUWghVgTCBkad/tcb9l4SrsOIMT2
sCqKbGbNeBGhzjMLao9vFIrqUrh3RqPT3qgmjvZji/1JMbGJ29OLJ7KwvOIREykK
CbTH0RuzFu0Py6IHIcAik6LH4ZMbUhZm4AWEnJ62Sbt+CtwHnAlFF/2mOfoksqBM
PZbDj8z15K9LHPLjdyArKsAu67O+bu7L8y8UFF2Fcb/+hRMtHKUV9SwICPQOWQFt
qy02qN4mjUivk2dzFvErR7+wNDgt9uSxhMqiAt3ewVYBhOqmag65TbAEHgbAINKo
K+a+w1eyurTCmjV3CXPpZzB8Qi5ATMRewL00yMxZgw5msU9U/e20LOKylz41X5Mf
kzQbvHHWQPTb+v7AZkt/C/xk2hjjr8YpphCXeXOtcMRrpI6fKncLeK+ig5QGqeaO
WoJvQzkQ7Lq7/ObkpSCLxp0SC9Rj0btCWNZllpbMfH6UOqBfciVcbHlZGBoMfv1V
eUA+NgtHVt9DxOps0c3u958pG+wOiVCSubkAFTNXY36q/jdMpdb2KxvgyqfJfqZb
rdHfjlwfTMhG3aLsLnObvLxAARrGHNtsTBHLh8mRhNVtHAxY8Iubf1IiaMvVsVt4
faPMumpa4E5FoSQ5v5a5mjyPe060SQxOBPJ9w7gzqmdYQXFIIIAootoovxhrx+bh
otrEU+BHarIpA4O4a3w/Vn8A/jgRM3hUT/n6zd4CtsPIdDqTepFcJ8WENGbZJ06t
lRngqLY2QF+4HNwn46LInn8UL+47oyTgbZPayqLAgNYL5zO+6qsad4dWKDOOYjcG
gFzUTuo7+cZHjQyBAOrLjuHigqIrotvvulRkCKe8fm3F2nUq1IwhnsFJMeRXF9pv
Lf21+605e0whlmPF5tRBAaXHLYSEp4GuiyQflzeJH2RNLZaOrRr2Op7XjvouAgHJ
pi7eA/M+dZI3RaFT5nn2OpqFosq/SM0KHF/Ci2CNI7K7zii8/ynvPhSh3eF5nv/I
Ug/m1pU0Ltci2SXapR6e0w3R1MiO4KLkihTaCr436Ew320BOPqYD7PpCZJ+yXjWa
eC8qaIe6tEfqxevPwb/Gca3UgvXyvSHyxSAcyE1Tz4Y0hdyOa3KA4qV9xJu0bbNE
LXfAoN0f5nmvULWuWTpEtiIdCpRkkAUqLEV8iu9ybCfwLY1Fs/s1vMncC5/7AQSt
l4Q1EjnEur5+TXFZgpawFObkZ+qrD1BaT00bvYWJ/OG0xCT8eD82OWap7FyrBh8I
+oQ5XDRsTOw8Z+h1Jmx5YikRZs9Z3TWOQoQBrep8nT2IldW0dtCICYFyWbJzN28e
MWF8RRFeOQVMM65z3yea3SvtkYWc1GJwF2H8lYAAeM7k8teWYCjAJqTh/GN6Z/4r
cMXjtPKGPRjQ5uh/bEEGCr+2IAXlIVm1kVkFG72VYwHGy2fyvQYv8sCMasOUmXzn
tfQSeiddl9c1PvHULkNHI79/3Zc223aWusn4FPZYfgSpwxcSZzGrKER04Re9Dtrd
xHUCZg5Mq4Sh70SdH1jcBfu06G2nU+yQc0eYAbQx1ZWp9etiDJ2Mo5dytx39KRe7
seYYzQ35y39NwVcTfh5hZvlh+cZnrZnMUD/P6SsXVR9M9AxRcPJx+w8DRgiJ+3gw
fjxrCayWF83i5epTB+DgMe4j1JKct2jaXQJJ3guEtlFTN3wHTH7/IpeJY8D1a3rb
eoq1Xui1R7cGS7vIBPyutxv8lriG6+F81Cxeyn5ns7FeVXQddF1CA423NdvVvT2X
lQSHHRYbJDeQodDw44vdrGuKmE0jv43yPt2InNGA748di0fDZCKV/lEcyTEQWfhW
4JoqQ3g+ebF+aEjiEWL0unRmhdAcwtdXJTZGQvr27ip7IqLZs2Ykl/xKeekKvCqf
40/EfCi5Wjd9nKGhIZRY9RjgXv/k4GcEY3elH2Dux7BrqQOBM1HpO3rwttTr6rZc
aXRGH4FtkBnsi46nXyrndkmWV8mZyXePbJT7OpsnP8ee4NiyaIaXBjJ9HyHIMt5W
ko//8Hs9diHy9twCecr2RmQotxxsVbSo4+93KnWYxNkhpL1Q1lNYBXurJMaH8ybY
ArceNaaQYcqIhwpujXnlEdD0e5caGy14lp5TLBSkOUCbO0/6XXXE18Rm4zZh4Y2Z
yuVYk08HqwLa3w77t9oKPDHA/hD3DCjyhi/aLZw2WRz4K3vK8iYzzlxZyl4dsM8g
e8wGwtUvFC4zaVmRGCVpqEgbwGOFUF0RFa0mesLAmj2FTOpMcBba2pLzaSK6Z0Ly
VrP+nno7f8DZVH4zbKGOqEOjiGhE3/L4jE9F1Helc/JOdV2Zzblcczm8+/NCBfId
bBCmT/KjVfSbxailzQTrREatuZ6nr1j4iLITe2TN2BA1AmNLgdMv+l9+cqR/5Gy+
2/Y8PtJtSK03jZNbjQzl25dmA8upQOiovrRnjXjbLXUUT2sFZgLx4uY/0aIm9nhR
a/xewYPRoadWX0hMT5vOy1FCS0AtvfS7OxlnR5Uylxz8d2Rb0hqMIHmOcZQ4f55U
WwnC1pDaebS57nRDyrJgVWULtuFCf6vfq87OWSJJwUSwgzd2sNl76tZHwh8Mntd6
SRc0dYcPqAQESQTwvqE8ItPeo7j3BXBCDgiqz5hGTKzN98oB6nfKSJnb+LDzRGoG
RRpaQYl61z8xVqic6mIM/TVgr2zBRcL3nXVr8QNfbTq6VUhLym5Y+O8SNsrAR3ei
4jNU7ios00+buRIdBDTlNDr4Zl+6ldfpdt2zip6dWiriXqJ1o0kJGx3QVzPY3K5J
MVtNXKuRcNG/m9vXN8Xuq5bclIN7c09h23Bhx/LWdOZG3EfA5cUSSA56vsHrNDK2
1gRuG9Zz5UoGJ5jK94y0fOwc64G40OdinXPZSsqO4LvL/yv7kB1FHoGF0gV/LyFY
vsFdMYU454RbVEna4eMpcCftqpuJrjt8ef0g/zlLDvgCGThjtbGsgmPyJ4agOVyI
rL8slmoQz1l9vdtNXVk6GAw2s62WFAPGrR5jJzFEWWZo+Yi/IiwuAcYNO43J4ysp
N1/YH+hVebs3lAibL9KM2OL3Kzu/LDa9YIdPyu+lgOh3B33awygIkvpb8R2CZy07
bnx5tjlXtfsjRwlcyV1mXXxI/8Ld8R7Q3LLlSzmsA764gFCQmqCqpg9AZ5Oknm72
akjCjKbGv+apfbIHU5O1B/JgrlR6IrOXB+OJpzMfYv0CBsdqckhObss7I9Eibjvv
yP1BcHLBj0Qyhc4C2RjFWjGvN7sud1iyUTGieaQXEyDU4ksiDeY7nHMIntinVGwT
9d9u+gV0v6lT7k26bO1VlyOPYAII60ZwUJ/c8L09OvReU88ZH3UuLMs2+ILEq1zq
kR4pIbU7EE/M5aG/RH/HxPmUKKLubxYITZoZ9NC7mpMatEQCFTk5idhXYQi9Xs2D
HJqBXG0hMAa1+6NUQSbsqNCVY/pHXvQGpAEoqyTyhDFprz4pP+4snaDWa54jrKrg
btgNDSaU/s26o2BREhhLqd3TZ6WFeXbWPHC7yA7R4TnAu8i8Yg0LKRZy0cbAGF/L
uCLk/bOFbO/7GMRp0JhEKcKiObzQzknDYIZNDtBGQw5pkcrWW/n5HNTM2Ts5eKvH
F9mJW6/8EaePdy6QturN8Y3AaNJ8EhCzcr30zEqOzG6/Sexr/85kreqltfXVUX3r
r9srQzJWOtXNLr3Y7ReEiXacF2q5+9tE+JbMdhtTZso8zp09RBn4zTrYHKwnCXA8
0D9vvRhpDg80vg8XxtDqrWb27eFhTuCKzgagGbOEcggHG40MbX46ptgRrcitaTRP
zdFvBGOSwUOQ2IH8jY06Qahrd/yRnr1l9hs9erfRhMqN8CmfbAarwMEuTqm1aU/S
WBBHqpCxsH97vL/6IcDltfCvOd6wrX7/AQYp2vxt30S8Eos4O+Ydts/AVzRgTvjm
/EKpeCzDTBYNWx3Boeb8cM+NciZWZmtgevgFxH+u+OxTNq/UzfFA/FByRw4vU41/
LKIYl51AkmMoEyW5/0znXJ+sH7m1+sIL1awg9YponmSy9cRvU2k3EXVAedSLkHwx
nYDst55Wb0CiIVHrK2k5o7Wwjosx7RMo8VFIHF5vUrEk7kpeOnEnu2NHcEqFKDHc
md+VoyQfCcoZrxblEJCKeFVzUuXWzQPsVn+pKmcMxKpotCGWcnPfhFJPS8GyOPKT
2VDJVV8DYBp+ZVev9UopIX2QgZk1br5Fl+0xGo64mScY3RffO/VKOx3K/b7ZpJcu
MqYz3tVmC6Sk6WRAx5q3D7x9jHr5M6VOfuEIEtEtxJlPGOyj///lKzHe4az2bSCJ
JEDE57iV2ixsTK1NbWaGFLm3OtM7FOGLW5fxMGlTp2t4aCbJsMc8ou4g2fx5e+6h
aJTPZ4tz/lYGpld4G101KELlnZO3Ss43CoSFZKRHL1jEZm+arC+ZPQR+DUJc5goI
iP/5hFfBhG3Ah/VwjPpxKDfRI8S8039gxw2X/icRGDyMOpdhId2JJbCl7MGDUPN1
oIxmaJJwkrmp0BgjVQh6GC5uFqZPQiZ3oRp9eu0X85qut+Km8TCcdMF1vI5ZTXoP
BJnibspKoftpy8e89r7tu4tywATTigCpgxjRSy/JAePYc/Y9vB7SyDxkY0hLFKrT
Y2JYZqVGp7vmh0bJ0nM7FdG+tTfiDDb7TnE6GGQR6YpNaf4cLF6d4kKovx2pmkXk
4YjPkyycy99Bfgz2IK2Kl7V3tAI9T71m0iPKK4rHB5Kbti1u3krmUEeuIY3w1AcD
Yu6ek0BrDcg1xdPmJXtjLm4UBkDzY2UAmqQDsHTBvmci8wPys0pMbtmjAcAzPaRm
DMQPzNFvtXOnQKTTnCJTBCIjMxME8d6DwSjwbyPv1FklkUx2WFIUFFbYW6eK4CGx
svJo0xOS2HtMABTKHB1mQvPXLpC2tH/Y9kcFDM48CUnRy2BMaZYwxx1ueyI5EQrQ
apKeHIFZQJ8qzh5uXkdJab3ZQ3itgZb8GiPSx6bzOXjBSZAqHHga4uay3dtzA+Z0
S3Ig67lLy/xiBnATOCEHhMqo5x08I27UaeudohIhAof8Z//0anzHOcXmqY7NthuY
JjkbrLchiKLGztKSmBDZda+wY3ydX4dJoF+FJeOq7TvL3wAz0MGMfhiyIqXvdMTZ
jQojE2Ok1gvFV2UWROAUL1KXy7Ejc0nnQvlDyyQQtSAwhsOCY88kfY6kXKT6e5ov
POstRgNcvQldDE4W1GO1xIkTPuTXO3PXy6O2OLIiY70wcPVZfx+ZnSHPFLo/Nj3c
Bt76RjRYYSeMX5rKzgogNNVLqbVy9hBTsipAPrMOU1NSbM6ljH3Co2fUiqGP/nak
fS9YhiZARkg6oiTg53WO++LCcR0TuHkj8GQZbtQEudrBr0R009NcoSeVsxMvTA37
PPp91tqqxnKjX9AC4Xj76xa45LZPSAg9tes09Mg8AbyQ6ajdZyntx/GNHrQ4lHMC
HyqJvkuuTJVZRYhQQ1AAAQaF1R2HYVMOuAKZKPGeI4gEnhzREg4HPo6iFtTND2oT
`protect END_PROTECTED
