`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0QvDr5c+3j6mGsZXXUqJ69Mx5TDeugcc7zpyOT1YpbKZN835tU894fgM+HZtl62
S/hjpsLoALe90y4ma368g1mbrnSvC95DTfRs8SpkzCY7P1TZprDzO1JQW5U0u1jc
J9riiONLVEYhuYq7PzoV1KY3A9riQ/bYaT826mt8s/mrJJaGolMTO7Yto9satXVJ
GARZFbJGRSs5fI1Orw4cL27fS9v6VXxIeXtIyWFdNSBw/Y1iugolWsdVevjB7tnT
bV68v5p25E53xmqqFPq9q+9qUThy0vySlBLfXpZP6xwBf8lqsDU+WNGyqigrQ/BC
1gt3nXAID3oWM0qHYpJW/O60bjbafJ65sTvvnxreQG+7gfWPoW8Bp75iYTJBRZSr
SMfu9evCeilJItS0sDu1B6egDQ5w9JdtFxkS2WD4OO6VibbHZDJftrTstyaph9sQ
O2SgpxiQBDW/fIqmhfBX1HciIDTD65qWktB4oVsr1vWdNfekng5+LlgQ229cpULD
jSSDEjn6HFcRjDOR99ODjH/ElLQBCJ/BN0zSUcJp727kPTFLvOvy4lu9PM0F4mRV
sgpSvq2vMdfd61OT9zrvHJbDqqDW/cPb7fP6TgbHZi/rWa03nMMrZ939Hc4C15rw
TI3mH+9/1LLwNs0QPF2lofF6P2NZVd6kKeDsjerl0PP9ozOf9jshE9Jq9T0YLsC6
eTyRjUFxzxFKZf90580Xr7H39RkbI2MlV/GO3l6dnn8MrK0Om5p4fLVuDxqb78s7
yuvDhY3GOmab0o7koUw1Q67no/xrr4bA6wb86X+GPWbP6lH81rSGYprx1b8Wweds
`protect END_PROTECTED
