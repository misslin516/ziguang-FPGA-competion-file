`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaMFxAlZZuv9dcv9lbKeT0sicGOBu8ITDGvvgCCTqrAaz8X+IH7TC/HgJ2/BAbSR
Xwlgik0x5LI0Q+6zmvY3n5gYOyF/r/dZOKEqM8Po3Sq1kB8QPVNyU0rLypNgFoWn
ul2Unv8ZMQT/2yjVse6JTa6bzLE8c4ieoNtKNL4doa5AIHbxQqvSSQesGH7ykjvT
yr+bXyPiB4h+F/1gS5IsPf5IUkdZEu0nTYgHYp3q4QWefenUKSzzypCDvVkTcIKa
lSBxKCSI0dq2R45RnnZ0ZBB6MyAt0WPfPDQaxMf4HsPJZQsbQCSEM0g3IDok0moT
auGkmmeUwvmxH4TURpHyC6TUcMlLDBMPHd/r0GR6XxouUDbNrO4KGCUuXYSiozs4
uW0JGp5yWi0Q/mAeqQpwIFcGggy0exqRHzoPr0VyZDK0mdZBw/poKhE8QNZTTjK2
KegvYns5lbcPecMVzHgSq7uzFLQk/hg/P7bYIs7VyoPwlx080AaNgpo+6zgHa/+/
rxl9kT2hf0/ojReFII1FkKaQpw89MH55TN/4yPf+yC2T29nlw4g9UKMFhrI7PrBD
fzvkhs1G0J3+NhwuHQmTyQHRHw9Oj+dndimmeYeeZwQbyxX4J0OqeShBQy7Ew4gJ
rZQnPMNPupX+kmeNh/doelc/8gyjuh4GHKwG3hTYfE9U2sNxZQRH3d1e0Qvb561x
BpIqQuumLBpaiicRV0Jp7HW4fES34YKw5ZvzWsJu6Bk3S3iWgEl/tjcnDC+X1IkS
ZM+YemCWCHnqZHESoEtV0dUw1zT5sGC8o3kkBkocQlm8l0mJMUlLGvOfAhUGh9we
1xNxQLgkbxyMxAxXPD7d68keyB90CuN8lDmCZYDLiQOcVAeQ9fwn/69SI4ztCh0c
z3OCmF/OEtZcghFzNAbrFhfw4GABvo0aYVBVsD0YAbdnsoSrby33RAanvi4IDdYY
Q4z8EfGRPVGoIt/v/H0kzxCsU8dwV9UjoHU5NjLU75n9oCgJTTssdRjRYlgFywtp
U6pIzErINrHJ38NeLQeHTlKMs6Yn9H9VvoNU5lDG4bmjxEsVlCkThAOuL9gi22UA
2+O1AibSAWbQ0vm4Fc+jAdU54/Khi6ybmmPXANVtW66jn5rtW64Jx9wBuqHDL2EW
QAvPTQ50o7u6i0+ugneypnNidr/EWo4XKG81tcUx4TQojCmCjBUejbFf6y2SMjXZ
ubaUjtDeP+5YyH0Q/L9qCQ==
`protect END_PROTECTED
