`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exskUmmwS/nhW6dWLSk4ZTn0tUYxwOngmo7WR3tzJZgwyhUD0dno9dymkUkk43zC
ogVwW77aIAjMmUEb2JIzd81sWuuowZ4kJKRc6ACXq0Bv34QrdYfrOTgrHa2arqNL
Q2UXoQLxnMrp80LHz/KQ/ZW6CF58QaiXPCONNUr/Ya8r6/uhGqa8hdD5EhK7eV2h
suGJwgichJc4jS7ppDocxKvVg+YzqRLjoWgtbO/jQOhBsrx8LOBfJWlSPVul07xW
MWeoqzVcQHF97V1C7O6pdQmnmzd/hqnm1hJk7tmeamDDu7DxoOU/PuJO/1it5iRo
v7IlDmFgAx09QTRr1gmhn+S4G0Et7i5ivzR+yYoj75z2pwdmYA0JxLH2gU5Xn2ui
Q1/KTwFzw3xp2R8WBJPXFsPd9F/hgD1peWSrWIgBG/DEASGXhrsBBH3knACEyTf+
9IitbqRQnaNDpkeMGWW5fVG/LUMMsMt8OzTiWHhssLOjdHCEuPox5fKzJD+xXypN
7TwTlsPq9ocvZCL6PMTurP8n1xYKhjGQLYjMeTgBGmSDB/OSCdb6iB1qLlJzOku4
VwQGfdvIMqbmjzceFtjcC9OVJYFI9WTPJgePISvm4zlyQ+i+AvQhBs5pBlMjDPIH
EMJjEzbXyQs0Zt7vdqAv7OzPpNGlUBg5CfmtmRSbqp/UokHiHNdEgETrMm8hcKWb
IFPoXYngYxHom6G3pPyiSbYj2N69EWVNnOQgHVWKSfGISG904UNdhrP3zL4+2c6Q
3rVmFm5pfSz+mpQvWyYAp2NUEdh0iC4i6tTskD+fRsvqlws9/9i7OISxvB8TLgPL
d1haL0A8nBzBdObBKdo22eMFHAPwdGc7VdvP35zzQRoHFlScwakXpXShWcCZKLjO
bGe2Oc9AkVBGU2+Gu76zOM9kr9WTyy89V54AWlQCi2Gjf8OvH+FZAcjOaC2vGlrk
W9UlxmO6huHc+HZYpahc4x/cmo10xFzXhfbezDU6XSz2X2EvsNwhdSsEn6H9xb2q
5ToUsHACqOQCZwqwXlOtFRiFhNmiQa0Ye0ZAcWYRtI2vRyCHaBUGN0PdjBuYnlS4
`protect END_PROTECTED
