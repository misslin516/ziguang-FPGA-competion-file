`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CfsWJ7srDXQhx/xIH93QxYQNKF/melrkLopjfQWrtS9qo4emgIiQpNuOPNgMhaII
jFGKRqm9B4Ui9UvYiOQbVclp0gerD+LsZoksgU+MN60mvAQcAcPhrjEhaliEl1M1
/jj39JEtKS9tJ//s9y07POPASNrRbb6S/Wbq1YQPxLh5vsMVxTbFC11pHELvFDKE
1xpVGvbvaLiLURuXvXOdOjNPgd6xpPmdbYVsrfKYnqKDpU0bDmwt56p3/rqOVe1Z
c7RpFLzVXNOHgleNjc0Bg5qYFYCkOWEpuMU4er1L74xvJg+s/EMuS1otvMNgsHJv
8HeRKSB8xgHA9gLGfHlEltfY+I8ZqLD3ZEf6cBHcVZaHDWoKxskWw0xOQoicTK4/
fHPj6HsLfCULghYySPnFHP7elvr+w7Gt2iVM6muORJXpuXpq7wz8RK9kAkyWBweX
+HcHco4E3MjDzsZcgC1eXW+dHadRzIIKk54YYK9EyzbkXmQhEtkcOPL19mO6rbjl
OPrrrf+E6fosUrFGfkeb5lBdgk7uSR4NzkVyibgSD+HV4RqmPnS7Mgi8UPszT+jc
88nVhTzxFWgZUCWrnObgBHQ/nRyAY2RXMwd5Gbvxz0c/tAMRwRTnDInhDy/EQ8YB
/5wEGCWdiFqbR3oaddTnx0SvgVrWW4LIXyhcgftI66DDP+07O3d4d5oCD1qUTGEr
ybI5M9qyUyxLv7tDy41FRX1gKZHszwCATj+7H4sVZiEQTCWHgDDxFQeGqozQJ1kq
CDAQkvj4v5xwiZb5/VpaFmickOLhAS9j17IGWPuYgeD/6ie0hDIrDrqCj/rg/H5e
ZymMyUuJnQGLuiWFEsSQYkkY645BlharDczigVzKNp6PxQDf/EPhgCC1Eh7LbCNs
yyHa84x5n1QTN28fUy72ZvhI/WgqgoLlhoX3uAfepCSQP1Z1u1h9nBgJTGALmeCS
icPKDQWdzXfPiuGmx3QuMf2DWMqvCu+SN9qO63D5As8NnL5zMRQo16qQl9JCa2kp
cROuw++cSn2pG+0pyyPxug==
`protect END_PROTECTED
