`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVUoWXwAQN/GwdU/f67nJ3LrWTYjUF4uQCDQat1tkbf3U40oeZ2Od090+hbRgGq4
e4SJWK6MGC6B8QRaHtyJiSqN3xgcX8/y2jMhm9D21AjS4ZweV5KDYrGGn5Q2pbHV
G16VwUqs25mFk13AAm4tYEzJRBpDrD1DSxGfskdbQ2WM6K7bpQBl7+ZwqkewKIDW
1yV2eXdZkrj9DzEfphwAlEDO0xHDGKegQ7nDRF0/CScYhbCy1HyoM+0IgVMHuhgK
hj2463kYGDIwecXw0ifSCReEXPU0yVp73XXQZx/mhL2MKLGgDcLkcLAwwpHn1Lq0
VmdDwsD+tLVuSUWEE402xZDr4ypanE5ElnYZ9lYMhoFhwWUN4ZLPxGBmBTFnOEzt
VT1D9ukYzQ/dyx5RYo636qXIhcdwqfRLJpDy1ltSX8rEKtpkly5Y0RKV7bbx419C
bxuv8QTTWZa/xsf5iK1oT3l/yDtyTUDIU2XWcVw7MJqLZGWrDurSGfr3OeF/+TwJ
qURCNOiCjr1/t4gxPy0kvIyTeVcOEmYj3MtrUiZOtPOrboIyICdIEhGCAWeIz6aD
voVb7RhD+NeF2BqYd3IADkaKmhYB1V4FRcv+66Qz5+jHXTdU78wjRy/ZtxNsSmiK
TQqbBznSilPZaD/Cf6a9zpg4jX6mcslXyj57QjFEWSz+Y77ViiUmeoVKgrlI7xC/
8d+r9TB7ZsOeEFNORhJIpN2tlRr+er47Fab4jnjequbuw8B9uEA5+Z1bOaa1WRAk
zwAgoH3mj+ijhN3kWE3xe9bxtp2AasbCWv9iQzvRcKz4zU163rpMfOnFkttE3Qqu
EzDit+j5jP4kAYCJxPX4Q1qyyzbUSjRR6DONMYbj2RZTtnUMB/jdwwdBPYOPT3nv
7wzHk2APHyF7jLB0Rl88+XjhM13JpbbXiCiZWoV0ONA67T6S1as/VroSLvLrvMDN
sF/KvOyF/MPGHoUBGZnH0BO0CxG3Qzr3PVMCr1fNjnd8y62thqAM+m/ibwmvR4pG
6iXymlEPuPNx1tZmnlsb7N4DjHgc5oI8UaViq3TVwusvIDZ6knVZbux9vZHm3ghO
21LGKCBhyax+XCw0je0BNsxmXkiZ1mqjVlaXDig+3nzwepbAgM7fdfId10jcZ+1f
mzMns2pgw73sn8rupOrR63E7DOKAzZSztp3uj1uL7/Dtf7H9o4FRrQQIaMJnzgN5
BpnBpNz/Fru4Xaqdu+4eWjsCDgOITdGyg6sJAPawjftPJGnt3ib0QQYf5Qx6IYOK
OnrufeIl/QBgXlPaCWlkQJMkuASkji6nvAafTydg29bmTvnytztSahtIhVUEFKff
XWctDEMa748nwdCm7lCVRTN3LGploMKKZ/XW0fT9do9lXubTC2Cn+f6hpxEZ8Yfg
LjSwrM/YeIuIUIxYtHWA7bEOhZH64PRShD8pVXK7SlVV8elp+p3m0pZxmvtCGbLB
u46XhpYhK4RUu+yuPuKY+OB/ospNyu32DTpgCQDEDVHItQ7HC0jRssRey6bJD+6/
XOUoxkMNO0WqJc01gOPHkP9RuvSPD89uO7TY02vw36hJs1AD++RkKQyZu5gN6ZVF
BXX4obg284O9LTZdGRupvp6067XY41Vy2fBl3WlsRB0a1z2XXLUMKd9Q/HDpfV+n
UN+QGjWnb1sUSFgBAOFYX/kmqvXcneT8RIHAQF5ZXTV02MnuvQcC9k0LwgoEZ184
9W1B2JUru+N52K/ftf0SQIl8j/BmlfqZAsJffJXDgvZdH3NbsrpBq+YQIOJ62X8+
n5+aoPMMe1Q98UB5PpEeFL2LrKtJpQtaIsdHYYSBO0OnJve9dYwF2uKVQ84mD48Y
/5NJsMOjRZxUyNrw+R0X9pBhbVX7acqnLWf9F/7cojL6hUgJ6jqwK701MrKjv73E
TtWYjYfmxpF4SRWOhKL+tv+WqLqyVA2g4/e+W0VvWUZ4tS2i722yinvGxZUD1x5n
MZVPe1gz6vy2XsMyeqCjdzFCGklLFX9lUa25xDdRLbR7rvRXPq21W/BRsCKbzP0L
dJmosdIPJOlVCQiOfjwJU2k0X6R9cKSx/HkTOgyXYaGFE/KC8ZzT4jHa4jzr/YJS
oChJMyWTB1kzlnA2dC26VPQxV4Df8D9e9RwhL5Vyv9NClNp74B8h1dL3hW2c/URi
oIZyT9DPEZ86pCF/GkEU0MTCP/RM37Rv9BKjLfYiiYB5vHhCWSyln+6XV1BtzKyt
GicNbeQLQe/36nCoDPIeLclFTpftLWo+gS8UGWszZurV0+apZ+pebuU9MH/xHXTs
geP0rn3FfC8nm2I5t3V17fsn+5yTvUWzJ683Vf/XSf+GCExkAuVl+4rN+TeySkWG
nmHEinP2czhZ3mAL9lMZRluijyFR9xJId96LX0bPm46KdzyBlUFB5C+ftkAMT/s4
Z+gpFQH6sYcPj7FA78pHHUrWqX1mmaoBOfQBp+Sy/4nt8XRKrJ9u16i6eJ/qqh4W
ZvqIgnKCo9hWcuBGVFgtfup7Gc0StJZ0QAMCujO5QTrGZr1AgERfYGehV3JQodRk
3MWGIIAqKSfMqHNx6qSSptFA59B4ENmogkxvGUZkROw=
`protect END_PROTECTED
