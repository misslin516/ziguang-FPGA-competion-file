`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvCPxLjpvOkWbO7hktZxeVf2cqRIjgPzS6KDP1Jxaxxkx6TP3m9zeduZs3Tz52hw
/nhbiw7Ny7y14OF9C8jDNPy9U1gYfLipo3fXILZ7BmWTJxa5Jegq1pVbjnYpLHNy
nQ52unLwYpSDhzVIK1YVbm9OsntRXmt9/JShLR+O3d7craVqpSp4f0uXO8o1aBak
VRf5ULocrVa0Vb1JfF0esLmjZqb71nnwb7aAiiaOXv8D2nGyQCtVuRINzZ0H4/gF
7Pl7pio+hZ9DI79FnsrScOC6bDi+CKsVoxkko84/zxDpH50FK0dy1FS/qtRxhtAK
7GrOH3HD8IkqpRXpdEckqfDWXlGeVzGcIykc4ux4pn5RdopOt8EqH0WFxQC/6GfA
DfG1NikCesgrSJbWR5UTgS5+KfULaiyp6mxM+gwRnmB31dGZqrnjNKIKCEkmi7Tu
Lhs3+DHMQ+S4Ba2qb7ahI6rPKG8BJRB+6pVdPJw/wCV+zAANpIuMMg93yCgqopw1
gQRrhX8pJIu2vsekhN6YOGv6VTgI9TOfVoNARDcWSwBtmuv55qZxKAgZZ4Za2un6
WFbXtoz6GktEwJK3anlxaI5dLS7pnFDk7Xpwj8Kr2K5Z1xb865ZoakQU7Zr/UGe6
fRoCgJvXEKwMjnWjJtMAOLxzHfuSDE0ze/fTwKV1P2ZNfdPI7iRF7V77Vo1fYnta
rxnLkeS2kgZcnfqF0p1xexrR+NKTc+STFn4ifU0kLH1SVydrjEwQ9WoKX1e4Mu6L
M+sbqVxLH0uHd3h1l4iHakV3yEJQAdvlcT0O2e4RZSw=
`protect END_PROTECTED
