`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
13cVq7u1MKBombftih0Y/WagMj+Yd12dsthSZnOcvsEh2Z25VZS+uyfG8c2GwXyG
Zyxe8So7ZpKlRx8vgXndNkYPdam66vObGJAuqmiY8quxufr2c0+8Ow+NEgHmK8k4
PoNSW7siR20t2I3yWVFSgnyJkphDg2KxcqW8drY22uHOnN4JCmGMf16y10/MI0Yv
o3/df+9x1i7Jc+zG2CbEKzgLV66mPtztn67IHQEe/h5SvHZmT4WFPqs+x0wvrfHU
xHV3uYAbzI12xnoap/A/Fy4pDtk3xAfEASQQ5lGS8xCHWcyyuux3lB9jjAYzwQ2N
QNL4vYd65/sNvRiIMQRhjb4t1aWrwWjpXyxIxxRa2QETtwJGYQHGeOWYH3Do3QNc
OFILjMWUne7jJTeqdDt0uGACmEcSjOx6d55CdxyP+fklU5wbOIP2/QZitHMufKWJ
Tgp7hXlibOIezKcg8Fp0NtStyT861SEu4sjLFSFRosmrC4X9HXOb46DY5tOaqa0W
Q3icLgeOyqfH7M4rYRxqwCJGiazZU65iZfmEjSOMc9UC4SHV38kw8wF7ZctvekvE
JecTa+QH60oCIs7hl1GqQg5fgn+fsC1QeV9AksMnjwhl8Yx6C1aCxMXbn+Cqv5wo
3laZnAfwOZID29869B6y7RRg7pCU9x8lrAWNG7rntA+W69QXnpMnVwjZ0OjIVCln
nDdIRDIDdi/1oesbhs40/01qfbP8pRIfQQFjXYmkUZnELiHFBquc+Sr9Tb0kD4oi
mDZnzPaCvzc4+joZPsYWq5nhGbgOLmQG+dwDdVMAoIf/anvSsE9nRS3kNeyNGCDs
X8CNbpFmIVXfDCc7lKSot01FNaWcKOPkhEONRuRSQl3engHUOvvTRpKK1GhIl/XC
/Ao35R/KMWPJoIeUNYNX5U2n5i7yfJzbyY1vHI7OFWxbrgTpI3tnjyb0yWxJsJMz
Z0CL1A8ON2K/k/qiDqBhXxL4R2rGZfdW7p1SGvQ1iYSuOXB/2J9mWm3J2Gi1oDLe
41Is+nDSTmTtjoQBoGSuB3ed3Es3QVEZT5ZLD9kYrhV1dtPoyUyPXf0ULgz81wfI
apSRnDlvdcTanFOo2zFYtqYh5MG0EyD0zqHiCYVXI58UHbu5j2yJi3kmNbkSXZvf
Se6lzHbOKe3etEic4kcX13TdljTyqk9xd3XDJybzVMHRmejmVmhh0uNSpAVS59Qg
nZNwjHoAMWMr22FjQEiuUxZFpw8yG5f/T+U2lIIoVwVN117BmbEjHfkvz8YqX15v
tw9Kbq1LxQyMjYmCMrmASdF9n46OAJAqFxAUeyRVYovW9gZ2QHxVeBLfcDdBUUNI
1sUZCsz35DA/v+srLljfxQ==
`protect END_PROTECTED
