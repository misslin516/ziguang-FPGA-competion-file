`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zGpR5XKXlAWyrGd0cGYICqOOlDbnDrUETjmsw3cjcYnKy5TXAGSeZ+rIA9UwbamP
ggUaRIruFdUGhGwrXQicWrlzqhYr/qrMoZRFGX9tN1wr8/D/4HL2nxnGcPCuoKb3
GHmxf5T8VtKnwp47pOSiYekahvFCaEIohBmRSoPkAjN6OA+xY/KxHI9Yjj+exC2z
gj772KiQ0j7VfoTNIjypCkcqy2JNUGWn7feu4LVMiqSSBAIySqKYvlaXVMfAuJ8o
2SlEuA1ixlFggiB7zYQ9PoyvurY0F1YVH6X9zZqPdNJF27rInFEAeNa60fyPevU+
Z5mYtT9q+BE11ASYWkJvRZfKzKUgMsdB7gPywBgW0etqs9DmtmnVDDCuVafAPdWi
yZSHmSk6xWiNvqCcs8bar02/UR4xcdEqnC1Sa4q32tLeBZcipx7qfUO8uTojPM1l
nh6pQODxdhhZxW2ZxFafnwmlRFln48Mz+lO7KfMavGhzSwj28FK4pr9DWedxhRxb
X0k0HgE8OoB66rFVy/eidxqFWOO5uEZflRDC/NY4yTmy24fbbcVUWLf/4wgjndCZ
hs2DtgxBWaFDCXdJG3AkRXuMrMJPtFK1gtVZ8v0nRuCyPYWdT8NYoX8GUUuf9gTl
2ltLeRJehCufA1AB4lX90stQEQvrVCc6T0PWJx11QIxCSKyUxOuJu9p3X9J+Wkub
WI+4znXORdkHSLTsj4DEcGThobnTo9Stkm+3XDv7rkM+qsaJb2CmDodE1MVRKI2P
VKtAqZQLz29aD3wvwA+gWovauzQOlz3ufGq9pxO+z6vSTY5MeVApG6MoNzD8EBUM
IgGDf9xvjNoES9pmeAHCym9xWoowlbsf7AyuXJgNIJovVKfVkDcrMhIEpugIxAeh
MdWBwZTbMwIe4bC1dpH1Z2wsExDZWAORjmj3HABR54EfkMg+/iadLNt+Io2CO4N1
nI7FCLalAE6SMiYi9l9gC87J4xz4y9XWpdTHWuV9Ct5OfC/hlBzl2tqt/ytgW34T
1KDkOyNg0XLpGSOa0/QlRSCiTeLEpX79kL+nBKRuAx0M6XkA8l2TSitGk3VxB6Rc
YgU9iz/5v4AqeUGzI7OVe2dymINPNm6EFUDcSy6wH19GrX9llvaLP0BsoZhPklHy
TK0lwOnhhUONnUnVIofeC0KLAgTilH7Pu+DHMNyjsSs8JK+W3++NzBiAQpUwjTVe
cG2sVI/fcFl9fHJ38a8Ifqep639fHq9ZbV2zAX7Qt2WAOn2CUroy2QaTABmFlKuU
U5nyroWN3AEJ76/VeaZmKA==
`protect END_PROTECTED
