library verilog;
use verilog.vl_types.all;
entity ddr_test_ddrphy_top is
    generic(
        T200US          : vl_logic_vector(15 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        T500US          : vl_logic_vector(15 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        MEM_TYPE        : string  := "DDR3";
        TMRD            : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        TMOD            : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        TZQINIT         : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TXPR            : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        TRP             : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        TRFC            : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        TRCD            : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        MEM_ADDR_WIDTH  : integer := 15;
        MEM_BANK_WIDTH  : integer := 3;
        MEM_DQ_WIDTH    : integer := 32;
        MEM_DM_WIDTH    : integer := 4;
        MEM_DQS_WIDTH   : integer := 4;
        REGION_NUM      : integer := 3;
        DM_GROUP_EN     : integer := 0
    );
    port(
        ref_clk         : in     vl_logic;
        ddr_rstn        : in     vl_logic;
        pll_lock        : in     vl_logic;
        ddrphy_ioclk_gate: out    vl_logic;
        ddrphy_pll_rst  : out    vl_logic;
        ddrphy_dqs_rst  : out    vl_logic;
        ddrphy_clkin    : in     vl_logic;
        ddrphy_ioclk    : in     vl_logic_vector(8 downto 0);
        ioclk_gate_clk  : in     vl_logic;
        ddrphy_gate_update_en: in     vl_logic;
        update_com_val_err_flag: out    vl_logic_vector;
        init_read_clk_ctrl: in     vl_logic_vector(1 downto 0);
        init_slip_step  : in     vl_logic_vector(3 downto 0);
        init_samp_position: in     vl_logic_vector(7 downto 0);
        force_read_clk_ctrl: in     vl_logic;
        dfi_address     : in     vl_logic_vector;
        dfi_bank        : in     vl_logic_vector;
        dfi_cs_n        : in     vl_logic_vector(3 downto 0);
        dfi_cas_n       : in     vl_logic_vector(3 downto 0);
        dfi_ras_n       : in     vl_logic_vector(3 downto 0);
        dfi_we_n        : in     vl_logic_vector(3 downto 0);
        dfi_cke         : in     vl_logic_vector(3 downto 0);
        dfi_odt         : in     vl_logic_vector(3 downto 0);
        dfi_wrdata_en   : in     vl_logic_vector(3 downto 0);
        dfi_wrdata      : in     vl_logic_vector;
        dfi_wrdata_mask : in     vl_logic_vector;
        dfi_rddata      : out    vl_logic_vector;
        dfi_rddata_valid: out    vl_logic;
        dfi_reset_n     : in     vl_logic;
        dfi_phyupd_req  : out    vl_logic;
        dfi_phyupd_ack  : in     vl_logic;
        dfi_init_complete: out    vl_logic;
        dfi_error       : out    vl_logic;
        rd_fake_stop    : in     vl_logic;
        mem_rst_n       : out    vl_logic;
        mem_ck          : out    vl_logic;
        mem_ck_n        : out    vl_logic;
        mem_cke         : out    vl_logic;
        mem_cs_n        : out    vl_logic;
        mem_ras_n       : out    vl_logic;
        mem_cas_n       : out    vl_logic;
        mem_we_n        : out    vl_logic;
        mem_odt         : out    vl_logic;
        mem_a           : out    vl_logic_vector;
        mem_ba          : out    vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        mem_dq          : inout  vl_logic_vector;
        mem_dm          : out    vl_logic_vector;
        debug_calib_ctrl: out    vl_logic_vector(21 downto 0);
        debug_data      : out    vl_logic_vector;
        debug_slice_state: out    vl_logic_vector;
        ck_dly_set_bin  : out    vl_logic_vector(7 downto 0);
        force_ck_dly_set_bin: in     vl_logic_vector(7 downto 0);
        force_ck_dly_en : in     vl_logic;
        dll_step        : out    vl_logic_vector(7 downto 0);
        dll_lock        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of T200US : constant is 2;
    attribute mti_svvh_generic_type of T500US : constant is 2;
    attribute mti_svvh_generic_type of MEM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of TMRD : constant is 2;
    attribute mti_svvh_generic_type of TMOD : constant is 2;
    attribute mti_svvh_generic_type of TZQINIT : constant is 2;
    attribute mti_svvh_generic_type of TXPR : constant is 2;
    attribute mti_svvh_generic_type of TRP : constant is 2;
    attribute mti_svvh_generic_type of TRFC : constant is 2;
    attribute mti_svvh_generic_type of TRCD : constant is 2;
    attribute mti_svvh_generic_type of MEM_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of REGION_NUM : constant is 1;
    attribute mti_svvh_generic_type of DM_GROUP_EN : constant is 1;
end ddr_test_ddrphy_top;
