library verilog;
use verilog.vl_types.all;
entity ddr_test is
    generic(
        DFI_CLK_PERIOD  : integer := 10000;
        MEM_ROW_WIDTH   : integer := 15;
        MEM_COLUMN_WIDTH: integer := 10;
        MEM_BANK_WIDTH  : integer := 3;
        MEM_DQ_WIDTH    : integer := 32;
        MEM_DM_WIDTH    : integer := 4;
        MEM_DQS_WIDTH   : integer := 4;
        REGION_NUM      : integer := 3;
        CTRL_ADDR_WIDTH : vl_notype
    );
    port(
        ref_clk         : in     vl_logic;
        resetn          : in     vl_logic;
        ddr_init_done   : out    vl_logic;
        ddrphy_clkin    : out    vl_logic;
        pll_lock        : out    vl_logic;
        axi_awaddr      : in     vl_logic_vector;
        axi_awuser_ap   : in     vl_logic;
        axi_awuser_id   : in     vl_logic_vector(3 downto 0);
        axi_awlen       : in     vl_logic_vector(3 downto 0);
        axi_awready     : out    vl_logic;
        axi_awvalid     : in     vl_logic;
        axi_wdata       : in     vl_logic_vector;
        axi_wstrb       : in     vl_logic_vector;
        axi_wready      : out    vl_logic;
        axi_wusero_id   : out    vl_logic_vector(3 downto 0);
        axi_wusero_last : out    vl_logic;
        axi_araddr      : in     vl_logic_vector;
        axi_aruser_ap   : in     vl_logic;
        axi_aruser_id   : in     vl_logic_vector(3 downto 0);
        axi_arlen       : in     vl_logic_vector(3 downto 0);
        axi_arready     : out    vl_logic;
        axi_arvalid     : in     vl_logic;
        axi_rdata       : out    vl_logic_vector;
        axi_rid         : out    vl_logic_vector(3 downto 0);
        axi_rlast       : out    vl_logic;
        axi_rvalid      : out    vl_logic;
        apb_clk         : in     vl_logic;
        apb_rst_n       : in     vl_logic;
        apb_sel         : in     vl_logic;
        apb_enable      : in     vl_logic;
        apb_addr        : in     vl_logic_vector(7 downto 0);
        apb_write       : in     vl_logic;
        apb_ready       : out    vl_logic;
        apb_wdata       : in     vl_logic_vector(15 downto 0);
        apb_rdata       : out    vl_logic_vector(15 downto 0);
        apb_int         : out    vl_logic;
        debug_data      : out    vl_logic_vector;
        debug_slice_state: out    vl_logic_vector;
        debug_calib_ctrl: out    vl_logic_vector(21 downto 0);
        ck_dly_set_bin  : out    vl_logic_vector(7 downto 0);
        force_ck_dly_en : in     vl_logic;
        force_ck_dly_set_bin: in     vl_logic_vector(7 downto 0);
        dll_step        : out    vl_logic_vector(7 downto 0);
        dll_lock        : out    vl_logic;
        init_read_clk_ctrl: in     vl_logic_vector(1 downto 0);
        init_slip_step  : in     vl_logic_vector(3 downto 0);
        force_read_clk_ctrl: in     vl_logic;
        ddrphy_gate_update_en: in     vl_logic;
        update_com_val_err_flag: out    vl_logic_vector;
        rd_fake_stop    : in     vl_logic;
        mem_rst_n       : out    vl_logic;
        mem_ck          : out    vl_logic;
        mem_ck_n        : out    vl_logic;
        mem_cke         : out    vl_logic;
        mem_cs_n        : out    vl_logic;
        mem_ras_n       : out    vl_logic;
        mem_cas_n       : out    vl_logic;
        mem_we_n        : out    vl_logic;
        mem_odt         : out    vl_logic;
        mem_a           : out    vl_logic_vector;
        mem_ba          : out    vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        mem_dq          : inout  vl_logic_vector;
        mem_dm          : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DFI_CLK_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MEM_ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_COLUMN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of REGION_NUM : constant is 1;
    attribute mti_svvh_generic_type of CTRL_ADDR_WIDTH : constant is 3;
end ddr_test;
