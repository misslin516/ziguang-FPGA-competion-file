`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFFQ+VAFEOAQsWXoq9VgzLLS/2dUr0oeHsInY/473+wML6/b+jqF5Fdycfx8AwYT
+MoHkU55ETIFVs5NGhvhh2hHIDWWJ+AHph/vOH8GHiYQ1M0R2OC142xzwZMCZ9UU
nVnpt57wX2gcFl2CU/nOSOZhhzK7DVbSjp/eAEP4fu5rVu7JJ/9uGWmSyRFSC4ax
JHqnmg88TzTMcqB7PHEylbQ5UT1B9HkZtyQfIJCf88mbFV4dhKmmcuvzvk/UQchk
kHjOmwHVW/ir99T6HPR7Q+d5+yNQ+QtBuLYRFJweMKNbq8wKxlswJRr87Gj3rpox
MeuJ39agWknt7dzUgH6F0zZGwluy0tY5f5/N2ubPEpqtMnb+kXDAq0hvZx6Q7BkG
KBlVqlTV7nzcIxsb3QCyElhxo4hqnR8QnQnfuI830SA0bOSOhXlFI85EuYXSsvOg
1+mHusI+UsAPgYT8vIdeoPl7RWe7NbXGGXVQhrqkfrlQEM6gcKTxcvCET52zivzZ
ZRL5OC8meaqIgsnuyWximNwJAe44CoC603uM/oltbwtzEbL9QTVGkHssY7kbrdeX
n0bDpiws5gooug5igy4GqrNn46tUOercDVlG7vDv7dhaMukyh99lERULEFhJAdy2
yF9QkEbMSPb/IlFBXZFRqUR8TRRRAjZkDfWOBGicV/4eQKLUlTJPfagt2ZzwHS3f
1ztSmoMsOx5o9i0ip1UzXXx5myYp9u+S6bqT7B9HDyGq33vDy7z2XtJv1HQVl7mK
bgX1aRiR/fh9hnAUqZ3lMtxGiEcreIOHkgOEnsRJygYNYIUuls76Zg8oM3N2nDe1
/O2Z89S7s8AAyA0O7nuXhVrOBB6ysY0CdaeIAo0mhJ8VfLDdPc/OsI9OKpKi4Aaj
QYppMXm2O7x44k1qhrtpFTBEn4K1STUELuny5FXtJZfUELehUEA6PPz3aQoQVRxs
ezTI4Ldif4HcconH90Amc9iO5wl3azidkDI5k+y9qbQ3emunTLRdmWFNmR/lM8Ey
IyRkVHoDhX/lwTF8sAEWLwHknxedRPNocQGIcjKcH0xjZKW4dl50ucvaSVtPQzYR
8CtzOQVoT3qhnh/mGt/R6SDsqlsmSt250s0xctSLt8c73j8RBiHLTmqgscCsy4Wl
eiQRwiEYQitybTPmPPH71JT20DAbD7yCPgKe+RERpKxAujxiIZWbC3KmCky32Keo
3PoFBfAIl7cCXPFi8qFb38DAYFYbV/1ZR6x03VRWX4EdPTRv3N2arqolNTL5ZWX2
cu2dtJT0re8rbASWa/BiFiax4J+qcni47jEFOufF1Emmwg+rtuU5iw06GfrIqqzM
w5mVYQc4wbdk/pQ9pXA1CDFMUnr7HaRpnFYwFLcdYJO74ueOCqvI082iWHzkQoqz
dq6GU21vja6IjWaXe9G7cV2scMCV44Q3qM+xgZ8XDSEci+qy2h+8oGWzQx5xl04S
UcEH3Salvd5h7xy0LGsyhtBwi/ipukQiqnAmg4JuItoHjNhfkW3nvQLpkWbyTS5G
7Fki7DI0LSzTPpeAiMV4kri+91QFJYp2oZRmTJcsEnVpwdm8rOM4H6eBe4Inloov
RQNslCrt1fVhgxVf9mGnxxwUE8ZiMtbkJmvuGBVNjQGaj+ZgnFH0cBVaoSxQzd0v
aPpC3snsG3UUXWDZq8bOibc+OneBYuJ4p+PCl8mOglwCsvrI6KpHyHzjFvn3RHnU
aIFSKlEVufkjFnNVEWpXGnMQdSOeHe5p0QfquBD+0/E2Lb//am15UkdEfPNB8cyL
shxBCNy+ZnjWNIiEbWdOPiGY96z0w5putcNorPd2g5aFIpameYBwE+jMniZKZheo
`protect END_PROTECTED
