`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6KLqId7a9kuTkTPnPwWksYwiTLeV6kKLSwfA38a2wMpBForY04Kq7ixGNUP4RYE
E/KLDj53STw7fSEI3YDhyARD2IqH9WIRyQxk5REfnI1/U241CjuuASp9OdYd07LD
QD88Ks1GUtLqp3sum7Xu32lqTj8dkEvUZsUv9Hbk5LpPrFGHwRR3AYXAIAmmpyej
n7vWCBQR50aM8vBvaT9VS+arYKLwK0V4mE414tA/yUM3ogG7/mgDpdTa5Y/hE4hp
M2772hbtB5HdCLEDAbUQb0kCu5NyRibhW1NA5zIKMKAybHBXAIVp+/CHClHh/dxk
2SCKIhU01zb0nHi3/w803vs1rTgwsUEiH1/eXVXu5d43ufqeTG0kzXr10dUBHizy
mEfcIq03KPNoERDhntlgWK1I3kGi+EkaAjM8VywZbkTOH7/BfLbc7iPj8jvCRo8R
9IvMJaFTnVxWRimCuozemvubFc7/UO7zeZAOZhv2PLsXaz74t8QMQI3eEbJL4soJ
bIk7rNJI05doPrhf6fQNUg6mF1tgcejt+xyG6GourUA86d7NUPvYPhtx9dKT+Kcf
joCpgEN0LkyFOefNB3+wWU8TocvaGnGc2DrbnBPdH5/NG9uxiT/raJ5Us+tqCJlU
KO/j8PyQ4zdPUqKRR4HVgLra29sXP0BvILexX42wYii/IS3V/SbjVeHXXq3pyYkF
oIlJlFRzY+wtqMIFU/XMaPtgxj/Y8UEtFLys06GfiOwtZCS+3wnVXITcP5Q1xv+p
pqycF45+ThiR7gSz9+3HJGPGpu3B0c7KmzyVbE4Zj0tXFDlN0aqH/ntfhVblBCVm
iMeonfOy/h3sX0oOm4g6N6XBqWia64G4CmaMfbdw7Waq9LeXUHEo9WUpnDV5Us71
MMOMmHo5Oi5fPb764PnweH3Ok8b6eI4zhopFhYbTspLFIRUBy81j/1Q7oOWME2Wj
OFjRi4qhGG7n2kyZ3e4k1ONCarhrPdC+MRzhG9UesD3Nm+7l2edEFd1h5aMkiJK3
vnCnM4epsOoYNczbArn4IRw8VMfgukgWUg8xR+95lclzQjgeMMGDb0Rqu4oxgw1L
ssiTKQ1xzQYEFsbjUSffC/QYIc7tGkNO/O7rap/ogBZT2f5o3Y8uO3HEPoC6FqD6
ysMLRQMvxnLFLHQzX0/dHQrWXGu2+TRDq8kqSagtp/eba8oZyDj9TedFe6jDWiEB
tePwb8I3pmxOKTaF/VmpHP6LmiGe4b7Q4uwTu59fqF56+NJJ+8zD1nvM0c7U/zUA
zv7LWuKplb/SXDcCzaIQk+xZY0R+XFWKZG/v+Pz2uTH6dQCE+C8shcWVoiQyd3Uo
0dnswnuR8Nq22JMTfAvbiG/vtYRo1ny8vkjEZKTqdXheSk2QqKEQ3P7L3J/KGB/h
FmCemeOMOUNmyFTdcbUIQqqooCoGdJdech+KOD3kscqD3JCrLysiRiS4hZiENoPg
0Auddeaxw0m6rOJnb/76KXnHPrIrfMitcreLNlN95ry481fLybNPg87a5bd8RlPe
EUeKajpbtuovOoQjXBMWoPN8GaEXAjMYkH+U5ur321nqY7KEsSPLN1npDErS99hn
sSlmjV+yagF5f1Uw29bdcx7pq8vdGUpfucBtDP4SovOX9QKn/up8B9nPyZKVUweJ
1j37LgZHaQW6p00wS2XhURUnL397wI5fbNC8h7y/w+UsKX8dfT9fEe7gpRkLOS7a
pYRme4CbYyrOi+uRIMgrHxhtuK3M/6SZUwfRCBas3e+7AQtSgtzBlRWl78Lu5Dsm
UbqqqXXRMh7ccryelnPenbvdw1kpgBO4yh5dIRlcKp0Wo8FmiuyLhQ0H6ZKdUsE4
L7SAdsqJGj5JH+ZhSq1JNYglgvqbBSR/VCIn4M7+2wez+5RGimaVfSsyC1S10/lC
zy4Fo3K8nAaC0muALkhhHhkDG+9gOaIUwV3LNGpwzTzlrA3v5GbQYFu64t6dc8vd
0TegpbPtXuGkQXIlBr9UKduf20isONKckW8KMZPsQ9O2FH1vJD2PtYtv9WiaYk59
1NSx0rr54F9yMQMerZhRnPK3bHpQsOawO0qNnTOKTooDGYDPpNndIrSpzgwMYysN
zOMLP30w759Hu0axTKAy9z08EB+WOiCY73sm6PWRPisL6JXBPpAKP4saadoJ8vts
XpAdclifuXY3X07ir2MG/CNFu6I3n7lvuxFEYn08jB8f8bYmRXFdAjJaxKYezn6l
ZXnClGv+JCVbrEEWCa4XQxIJSTgoHoGeDZDyH+BU6vIhWvW2Lf/I423yIIuu6rbd
UDETcpySGH3rXrjJ8+1Kfa7MOit4uCfcYCMA5TZeC3tZLSc37IKJtlOSQNESlM4C
XplpYWvlbWsd0s19Z64lho9YXLGx43zhX+bEkPYCf+ytd+J6z8exeDEYeOx1Vkss
YE01cz7z+1YcIOp8AOOFxyV7wkjHXlT+4l2t/EtxkPEmCix9MHmuxFShsQFuuvln
tCV6EhL131XuYNvx21ntICrWF6mt/1AqyyeLtUCMXX78yj8X7PrdRlBLL7IAozrL
VDajV+9pNLbE/DBD4po6bukM18cZVYXAd0wYsc0n/Kc/hx8KrtW3BIFucsfHKNEL
4n82VLzoe/dGn5s7gtzNk3pzHsgVGMPS/ZKWngphHYF4wdDWiBi54JVYV3PHkXh7
EkJRuO3JCwF2KWMDLlDF/UKk+VCgHRj7PjYuugDHz8ncTbFxRiprgqgnVqWSD5yW
QCmOjg+CKw1v5kGzezO+XYfEVU0Y4k2JgZU63UC5/8lS2H229J1bfw/S4xgGKoHK
uahbIc3DgcTGd3PPAjZAtHFNahTis6ke1MnZENXPpEyBu3bdn9OmvGMrpvTemvJY
ey0WtN3ufNEarpetxfkaetyAsaaRP3D7EvuxAZJXlLd0F75uh/V5ARkN9zdKemcw
XloN7bej11ahlC2F6xEZYSj3BeCb/Ymwpja/p7v8tloR4McqEG0dZwD0G3s+IZX+
R4ZcuQ3wXX53MxXxEXl3ZW5Iwcal/Q0kVP9tO+3377tcBOY6JJ2X+40/XcWFwomM
a4r7wVEFQ8NAc1vIPU1HuuoR/OAShPEi+OMxyYyyp/ypM1p4HNbndrnGVsiplR1U
NrGUEgGDFGwAl+qHfiTDWsyk0MfT3fva4zujs+r9psY=
`protect END_PROTECTED
