library verilog;
use verilog.vl_types.all;
entity axi_bist_top_v1_0 is
    generic(
        DATA_MASK_EN    : integer := 0;
        CTRL_ADDR_WIDTH : integer := 28;
        MEM_DQ_WIDTH    : integer := 16;
        MEM_SPACE_AW    : integer := 18;
        DATA_PATTERN0   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        DATA_PATTERN1   : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        DATA_PATTERN2   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        DATA_PATTERN3   : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DATA_PATTERN4   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        DATA_PATTERN5   : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        DATA_PATTERN6   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        DATA_PATTERN7   : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        core_clk        : in     vl_logic;
        core_clk_rst_n  : in     vl_logic;
        wr_mode         : in     vl_logic_vector(1 downto 0);
        data_mode       : in     vl_logic_vector(1 downto 0);
        len_random_en   : in     vl_logic;
        fix_axi_len     : in     vl_logic_vector(3 downto 0);
        bist_stop       : in     vl_logic;
        ddrc_init_done  : in     vl_logic;
        read_repeat_num : in     vl_logic_vector(3 downto 0);
        data_order      : in     vl_logic;
        dq_inversion    : in     vl_logic_vector(7 downto 0);
        insert_err      : in     vl_logic;
        manu_clear      : in     vl_logic;
        bist_run_led    : out    vl_logic;
        test_main_state : out    vl_logic_vector(3 downto 0);
        axi_awaddr      : out    vl_logic_vector;
        axi_awuser_ap   : out    vl_logic;
        axi_awuser_id   : out    vl_logic_vector(3 downto 0);
        axi_awlen       : out    vl_logic_vector(3 downto 0);
        axi_awready     : in     vl_logic;
        axi_awvalid     : out    vl_logic;
        axi_wdata       : out    vl_logic_vector;
        axi_wstrb       : out    vl_logic_vector;
        axi_wready      : in     vl_logic;
        test_wr_state   : out    vl_logic_vector(2 downto 0);
        axi_araddr      : out    vl_logic_vector;
        axi_aruser_ap   : out    vl_logic;
        axi_aruser_id   : out    vl_logic_vector(3 downto 0);
        axi_arlen       : out    vl_logic_vector(3 downto 0);
        axi_arready     : in     vl_logic;
        axi_arvalid     : out    vl_logic;
        axi_rdata       : in     vl_logic_vector;
        axi_rvalid      : in     vl_logic;
        err_cnt         : out    vl_logic_vector(7 downto 0);
        err_flag_led    : out    vl_logic;
        err_data_out    : out    vl_logic_vector;
        err_flag_out    : out    vl_logic_vector;
        exp_data_out    : out    vl_logic_vector;
        next_err_flag   : out    vl_logic;
        result_bit_out  : out    vl_logic_vector(15 downto 0);
        test_rd_state   : out    vl_logic_vector(2 downto 0);
        next_err_data   : out    vl_logic_vector;
        err_data_pre    : out    vl_logic_vector;
        err_data_aft    : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DATA_MASK_EN : constant is 1;
    attribute mti_svvh_generic_type of CTRL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_SPACE_AW : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN0 : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN1 : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN2 : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN3 : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN4 : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN5 : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN6 : constant is 1;
    attribute mti_svvh_generic_type of DATA_PATTERN7 : constant is 1;
end axi_bist_top_v1_0;
