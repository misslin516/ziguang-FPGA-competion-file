`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnN2HZL5YEp5GvPdry3HKGvyE0eQjo9mf806MGpYypbrT/WGQ92ceuuvDHcQ3rBj
36RyVJoe9D3EUp8xwUHs/LhdiVl9pQEMo9vVxwbUh6UTGLYROs9lefGJQc5isfQ6
No8nK958R51twnS8nIMLu6FxhdREmbwUZYi2oL8Ndowoe9/WVT37aQyWRv9qXF88
BHPG9MTtWD9gE3SMXiposPwWAz/amVOARr5mhaRKpAW1DF4AJoYsq+yw9J+QRYQ0
+JbV6pNa5m47JZRUSLSo3nE8velruCaXdWySYzZSoOEExs8OM+QeTD85T99teaim
lkgCzYaPZi84lllwrCD00sUJGiDJ7sa5wXwkoFEgqWmWhSggp0rFrjgx2GC0pcCU
pW9LdSJVD+aS6i76/LJOjbmGikysM2boE7Ivqur18BF6KWWbZo6NcGxR+kU1JheZ
lf/94g9gBYMMPEpYBqhOMAh/emBZXlAOqHPjM9qPUJ6+Ki6ZhE5k8JANp9tFIYE4
Vb4+SJCKUtsxgenGNFKYmMk22hpPGM7PiyFs+6InDnrN4/vH0Ws6olTTyDDfI+3e
AVa+z2Oxjx6aURmtlLrktrL06YUJ++hXzzXdHzPYmJSzEovSpGWNaqA660144Xa7
85MdCkIcJr4dLslyyvG+nkMDgmZJt/VRsvTOYkNeTF1aXgb61nNd/gOWByNgtZa9
hlSuwZ0UbT+CMrbS5nEuZHViZybi0ZqDSXGjY6aFTRLy9jp9kQLrBF3UiLg76y5L
Ew0rSfdhyKoVT01wg1B93OK0ot8i3WVG0OH40w8D0azp8CrTBMYVb+w0Yv//RdwC
sHHgph5zhuPmsgekxqQAEvxo6CaYeID6/RkTeUzlFilArNTOx0jMvcTHx/cBDEWj
l8YQXiPiDH5yM9x32LZRJJpaRnmlmheRtbsY2XKE3PkYNqCC44rJqCA9hT/8nRJP
CZfrne21Vosm+jA6e1ng5ginzmrPD7hNn6qWoq9izZC6n37HPEzam3yyVOqD2V1A
h1ykGHYI00XorHFVjseXOizSk7YtiGt2oKES4fgWkYSWaWDiQtp3I0B9geZW4Dhs
vxCYrWQHh15UOJqcBFIB+t+mjLilfoLrgIKhCqC+sJT3yj/cK8rEpPCUE1j7AD72
CBuQ1LeLOVkJM/Umbggfn6CZvO1qMbm1scXko8NkX52sVLc2+6OG0vxnwfHvWPSY
r+hlSIrQeexEwzGRJQ89/5cdEr+2jqsExOoz4WzLvyhWKEA5z2VuEH8QkNsMMeug
dPxoxp0cS8F0XOgCZOevlLfKxRv4gOHCRfrOG9+NSfJjzPTgt8RCFpNSW2GgQch+
jwdc2xPLRue3Bm+NSEzgPFnXjRUnTvaYKhkYmVZLlZsrK4YDqKqcOaqJF4yLlvYL
Sg6MnvS4MhRFrDEffNdQMRm9+FHRODLUxIa1tiEr97251F1u9/xr8xdtP/TijX37
Uoct43CJGd4qoYbwmsP98+qCg4rk68cbOFxDs7z0sU72tFhFMsHr6xQziuQAoVLB
hsplWyAS3VsBKDddXOlHFtccmsd5ly34GbsDhKu2OD7F6O0HyVrqLhZIzVIcjNzZ
Ny+P0+bK6CPavhLbVh1eP2xwMB0jS2duW94DtI2O1g/SqafJ3vewecojVsF/uCLZ
agO8VgvuT3Qn87zl8eC2wrRJHCCPULChit9owJBSoC1xKpQD949bQJ0L8+/3heDW
VKBBRPG+YtL/Ol3KQJPuPCh8F26YmwZu9PELW6p+sPkcoxLFllnW8LUjcQkgD3Bo
yNODRtdrh+dM0c2c7fY5Du3r6PLkEjfE1U8pI1RbaBXOgJK9lARhdGWD6FeWRmGf
p63fhJ8Mk9VBZEjfDm1mxSGW5vfQykY85xUPNzUR5l9VR5YA+eGPfOY/5ZIaf+Eg
d5USm6mtRhx/FUss9K/DNnsUvQlb4sOifOYTSvh2JvGaetkrwMFr/860qInn+dYd
y7wW7NJeiI88/hIl9oyvbOQ+PPaU2Q1CDf6rov1DB2QdMT71IVyDbuEtQxVNGe2t
hRyPWD3drR3S/s6sueq9o6kxmv6KO/RtlLJWR3iismWUkDfZml80u/ee7qAGz4CE
JjK+Rt7bhwZmOYtXlqdIv9BwAQW2HGP0sXNYV99YMkONxKBnW3eL+32iYmrjMbVg
R1G7O1tGmMUp649Egty20ebDOplm7SEo9vfGN9/PYOsMrZfS5Qrc3E2a9IKrsvUV
M6dKO/VoTW+DivbvnezNqxYmPqDD74Gna2Gk6e9U+qVXotGRXzlaQsvAAtMXDGGf
ELUpBFy0J1KIPnyngA7hKqYiJqJLrrDy4O00eQJBMWZtZMO/qmVQSFw2+kmv3IJ2
ZcF5MTKy8qaE8k6VcbhVX7sMz/3OSP5D2giM7exNFaVnP56ThwjezSubbgcC4+sV
cJcDLM0Q+L/8rPZXsrwgq2JTedc11NcyQIsr7DhH170c0xS8Z1IXtbCD823PUfvR
05gNgvFmrqHpbag/gcg4NqfFC42eO892jVJqfmlr1LOeMrdliAFUc2xWZGdsmDUv
62vSPa3JYAGP8FmnolbZvYL80TdYYKX+0dKczn/9qqCcujN7avqX1ZOpYmcSUkNT
Zl5MQFBQaLT5R7LMDAOBI4t2TJ/h85RtT3WgMYgTmGcY9wneaaxDQzlsOyAcmPe4
3qDnFUxUy/vGHEEWxPZhhRrxI6c+pECGLqqyX11Ob80JU8INKyvabyI1nVcaeQrW
5RwjxcrfU6naad6TPlbUB1ocAhHyxM8wQ85AHyRoqpZ5UT3EwqhY2sK2dew9fXN6
`protect END_PROTECTED
